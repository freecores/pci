// Xilinx Verilog produced by program ngd2ver D.27
// Command: -w pci_crta.nga crta_time_sim.v 
// Options: -w -log ngd2ver.log -ti uut 
// Date: Thu Sep 27 04:18:22 2001 
// Input file: pci_crta.nga
// Output file: crta_time_sim.v
// Tmp file: C:/WINNT/TEMP/xil_23
// Design name: TOP
// Xilinx: C:/Foundation
// # of Modules: 1
// Device: 2s150pq208-5

// The output of ngd2ver is a simulation model. This file cannot be synthesized,
// or used in any other manner other than simulation. This netlist uses simulation
// primitives which may not represent the true implementation of the device, however
// the netlist is functionally correct. Do not modify this file.

`timescale 1 ns/1 ps

  module TOP (
    RST, IDSEL, STOP, FRAME, PERR, IRDY, SERR, PAR, TRDY, DEVSEL, GNT, HSYNC, 
    REQ, VSYNC, LED, CLK, CRT_CLK, AD, CBE, RGB
  );
    input RST;
    input IDSEL;
    inout STOP;
    inout FRAME;
    inout PERR;
    inout IRDY;
    output SERR;
    inout PAR;
    inout TRDY;
    inout DEVSEL;
    input GNT;
    output HSYNC;
    output REQ;
    output VSYNC;
    output LED;
    input CLK;
    input CRT_CLK;
    inout [31:0] AD;
    inout [3:0] CBE;
    output [15:4] RGB;
    wire XON;
    wire \bridge/configuration/C343/N5 ;
    wire CLK_BUFGPed;
    wire \bridge/pci_target_unit/pci_target_sm/S_345/cell0 ;
    wire N_RST;
    wire \bridge/configuration/delete_pci_err_cs_bit10 ;
    wire \bridge/configuration/C390/N3 ;
    wire \bridge/configuration/delete_pci_err_cs_bit8 ;
    wire \bridge/output_backup/data_load ;
    wire \bridge/out_bckp_tar_ad_en_out ;
    wire syn17116;
    wire syn179878;
    wire syn179881;
    wire syn20486;
    wire syn20502;
    wire syn179882;
    wire syn179883;
    wire \bridge/output_backup/C3/N6 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C155 ;
    wire syn179894;
    wire syn20532;
    wire syn20538;
    wire \bridge/output_backup/C3/N12 ;
    wire N12384;
    wire N12360;
    wire syn177396;
    wire syn177397;
    wire syn179931;
    wire syn20564;
    wire syn20571;
    wire syn179960;
    wire \bridge/output_backup/C3/N18 ;
    wire \bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ;
    wire \bridge/pci_target_unit/wishbone_master/N3069 ;
    wire \bridge/pci_target_unit/wishbone_master/reset_rty_cnt ;
    wire syn19555;
    wire \bridge/pci_target_unit/wishbone_master/N3068 ;
    wire syn17106;
    wire syn20598;
    wire syn20611;
    wire syn180003;
    wire syn180250;
    wire \bridge/output_backup/C3/N24 ;
    wire N12545;
    wire \bridge/in_reg_frame_out ;
    wire \bridge/pci_target_unit/pci_target_sm/S_291/cell0 ;
    wire syn19671;
    wire \bridge/pci_target_unit/pci_target_if/norm_prf_en ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_control_out[0] ;
    wire \bridge/pci_target_unit/del_sync_burst_out ;
    wire syn24500;
    wire syn180012;
    wire syn20635;
    wire syn20641;
    wire \bridge/output_backup/C3/N30 ;
    wire \bridge/pci_target_unit/wishbone_master/N3071 ;
    wire \bridge/pci_target_unit/wishbone_master/N3070 ;
    wire syn136384;
    wire syn136386;
    wire syn20662;
    wire syn20672;
    wire syn180067;
    wire \bridge/output_backup/C3/N36 ;
    wire syn20688;
    wire syn20701;
    wire syn180098;
    wire \bridge/output_backup/C3/N42 ;
    wire \bridge/pci_target_unit/wishbone_master/N3073 ;
    wire \bridge/pci_target_unit/wishbone_master/N3072 ;
    wire N12478;
    wire \bridge/pci_target_unit/wishbone_master/N2993 ;
    wire syn16933;
    wire \bridge/pci_target_unit/wishbone_master/C81/N3 ;
    wire syn16925;
    wire syn182174;
    wire syn180107;
    wire syn20720;
    wire syn20726;
    wire \bridge/output_backup/C3/N48 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ;
    wire \bridge/pci_target_unit/wishbone_master/N2994 ;
    wire syn182179;
    wire \bridge/pciu_err_addr_out[11] ;
    wire syn20737;
    wire syn20738;
    wire syn180176;
    wire syn180183;
    wire syn20759;
    wire syn180180;
    wire syn180181;
    wire syn180185;
    wire \bridge/output_backup/C3/N54 ;
    wire \bridge/pci_target_unit/wishbone_master/N3075 ;
    wire \bridge/pci_target_unit/wishbone_master/N3074 ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/map ;
    wire \bridge/pci_target_unit/wishbone_master/N3003 ;
    wire syn182224;
    wire \bridge/pciu_err_addr_out[20] ;
    wire \bridge/pci_target_unit/wishbone_master/N2995 ;
    wire syn182184;
    wire \bridge/pciu_err_addr_out[12] ;
    wire syn180219;
    wire syn20788;
    wire syn137911;
    wire syn180212;
    wire syn180222;
    wire \bridge/output_backup/C3/N60 ;
    wire \bridge/pci_target_unit/wishbone_master/N3004 ;
    wire syn182229;
    wire \bridge/pciu_err_addr_out[21] ;
    wire \bridge/pci_target_unit/wishbone_master/N2996 ;
    wire syn182189;
    wire \bridge/pciu_err_addr_out[13] ;
    wire \bridge/pci_target_unit/wishbone_master/N3013 ;
    wire syn182274;
    wire \bridge/pciu_err_addr_out[30] ;
    wire \bridge/pci_target_unit/wishbone_master/N3005 ;
    wire syn182234;
    wire \bridge/pciu_err_addr_out[22] ;
    wire \bridge/pci_target_unit/wishbone_master/N2997 ;
    wire syn182194;
    wire \bridge/pciu_err_addr_out[14] ;
    wire \bridge/pci_target_unit/wishbone_master/N3014 ;
    wire syn182279;
    wire \bridge/pciu_err_addr_out[31] ;
    wire \bridge/pci_target_unit/wishbone_master/N3006 ;
    wire syn182239;
    wire \bridge/pciu_err_addr_out[23] ;
    wire \bridge/pci_target_unit/wishbone_master/N2998 ;
    wire syn182199;
    wire \bridge/pciu_err_addr_out[15] ;
    wire \bridge/pci_target_unit/wishbone_master/N3007 ;
    wire syn182244;
    wire \bridge/pciu_err_addr_out[24] ;
    wire \bridge/pci_target_unit/wishbone_master/N2999 ;
    wire syn182204;
    wire \bridge/pciu_err_addr_out[16] ;
    wire \bridge/pci_target_unit/wishbone_master/N3008 ;
    wire syn182249;
    wire \bridge/pciu_err_addr_out[25] ;
    wire \bridge/pci_target_unit/wishbone_master/N3000 ;
    wire syn182209;
    wire \bridge/pciu_err_addr_out[17] ;
    wire \bridge/pci_target_unit/wishbone_master/N3009 ;
    wire syn182254;
    wire \bridge/pciu_err_addr_out[26] ;
    wire \bridge/pci_target_unit/wishbone_master/N3001 ;
    wire syn182214;
    wire \bridge/pciu_err_addr_out[18] ;
    wire N_TRDY;
    wire N_STOP;
    wire N_DEVSEL;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N147 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/S_13/cell0 ;
    wire \bridge/pci_target_unit/pci_target_sm/stop_w ;
    wire \bridge/pci_target_unit/pci_target_sm/stop_w_frm ;
    wire N_FRAME;
    wire \bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy ;
    wire N_IRDY;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_stop_critical/syn67 ;
    wire N12476;
    wire \bridge/out_bckp_stop_out ;
    wire \bridge/pci_target_unit/wishbone_master/N3010 ;
    wire syn182259;
    wire \bridge/pciu_err_addr_out[27] ;
    wire \bridge/pci_target_unit/wishbone_master/N3002 ;
    wire syn182219;
    wire \bridge/pciu_err_addr_out[19] ;
    wire \bridge/pci_target_unit/wishbone_master/N3011 ;
    wire syn182264;
    wire \bridge/pciu_err_addr_out[28] ;
    wire \bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg ;
    wire syn182641;
    wire syn182642;
    wire N12616;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0 ;
    wire syn23757;
    wire \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr ;
    wire \bridge/pci_target_unit/fifos_pciw_full_out ;
    wire \bridge/pci_target_unit/wishbone_master/N3012 ;
    wire syn182269;
    wire \bridge/pciu_err_addr_out[29] ;
    wire N12351;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2619 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2618 ;
    wire \bridge/pci_target_unit/fifos/pciw_rallow ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2621 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2620 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2623 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2622 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2625 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2624 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/err_recovery ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/write_req_int ;
    wire syn60010;
    wire \bridge/wishbone_slave_unit/pcim_if_rdy_out ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ;
    wire \bridge/pci_target_unit/pcit_sm_addr_phase_out ;
    wire \bridge/pci_target_unit/pcit_if_read_processing_out ;
    wire \bridge/pci_target_unit/pcit_if_norm_access_to_config_out ;
    wire syn19927;
    wire \bridge/pci_target_unit/del_sync/req_comp_pending ;
    wire \bridge/pci_target_unit/pci_target_sm/wr_progress ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_request ;
    wire \bridge/pci_target_unit/fifos/pcir_rallow ;
    wire \bridge/pci_target_unit/fifos/pcir_clear ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/change_state ;
    wire N12359;
    wire \bridge/in_reg_irdy_out ;
    wire N_GNT;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C262 ;
    wire syn18858;
    wire syn18863;
    wire syn18937;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/C355/C3/C1 ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/C333/C3/C1 ;
    wire syn23402;
    wire syn18958;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/C311/C3/C1 ;
    wire \bridge/out_bckp_frame_out ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C4/N9 ;
    wire \bridge/pci_target_unit/fifos/in_count_en ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2 ;
    wire syn18899;
    wire \bridge/pci_target_unit/pci_target_sm/config_access ;
    wire \bridge/pci_target_unit/pci_target_if/decoder1/S_37/cell0 ;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn51 ;
    wire \bridge/pci_target_unit/fifos/pcir_wallow ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0 ;
    wire syn23568;
    wire syn182579;
    wire \bridge/pci_target_unit/fifos_pcir_full_out ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/almost_full ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/data_source ;
    wire \bridge/pci_target_unit/del_sync/N1246 ;
    wire syn23138;
    wire \bridge/pci_target_unit/del_sync/N1245 ;
    wire \bridge/wishbone_slave_unit/del_sync/N151 ;
    wire syn22149;
    wire \bridge/wishbone_slave_unit/del_sync/N150 ;
    wire \bridge/pci_target_unit/del_sync/N1248 ;
    wire \bridge/pci_target_unit/del_sync/N1247 ;
    wire N12467;
    wire syn182004;
    wire syn182005;
    wire syn182015;
    wire syn182018;
    wire syn182016;
    wire syn182017;
    wire syn182021;
    wire \bridge/pci_target_unit/pci_target_sm/same_read_reg ;
    wire \bridge/pci_target_unit/pci_target_if/same_read_reg ;
    wire \bridge/wishbone_slave_unit/del_sync/N153 ;
    wire \bridge/wishbone_slave_unit/del_sync/N152 ;
    wire \bridge/pci_target_unit/del_sync/N1250 ;
    wire \bridge/pci_target_unit/del_sync/N1249 ;
    wire \bridge/wishbone_slave_unit/del_sync/N155 ;
    wire \bridge/wishbone_slave_unit/del_sync/N154 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg ;
    wire \bridge/pci_target_unit/wishbone_master/C981 ;
    wire N12119;
    wire \bridge/pci_target_unit/wishbone_master/C960 ;
    wire N12118;
    wire \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp ;
    wire ERR_I;
    wire \bridge/pci_target_unit/del_sync/N1236 ;
    wire \bridge/pci_target_unit/del_sync/N1251 ;
    wire \bridge/wishbone_slave_unit/del_sync/N141 ;
    wire \bridge/wishbone_slave_unit/del_sync/N156 ;
    wire \bridge/pci_target_unit/wishbone_master/N2983 ;
    wire syn182122;
    wire \bridge/pciu_err_addr_out[0] ;
    wire N_IDSEL;
    wire \bridge/conf_pci_master_enable_out ;
    wire syn17745;
    wire syn24559;
    wire \bridge/conf_wb_err_pending_out ;
    wire syn178469;
    wire \bridge/in_reg_idsel_out ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/lock ;
    wire \bridge/pci_target_unit/wishbone_master/N2984 ;
    wire syn182129;
    wire \bridge/pciu_err_addr_out[1] ;
    wire \bridge/pci_target_unit/wishbone_master/N2985 ;
    wire syn182134;
    wire N12311;
    wire N12519;
    wire \bridge/pci_target_unit/wishbone_master/N2986 ;
    wire syn182139;
    wire N12120;
    wire \bridge/pci_target_unit/wishbone_master/N2987 ;
    wire syn182144;
    wire \bridge/pci_target_unit/wishbone_master/N2988 ;
    wire syn182149;
    wire \bridge/pci_target_unit/wishbone_master/N2989 ;
    wire syn182154;
    wire \bridge/pci_target_unit/wishbone_master/N2990 ;
    wire syn182159;
    wire \bridge/pci_target_unit/wishbone_master/N2991 ;
    wire syn182164;
    wire N12520;
    wire N12521;
    wire \bridge/pci_target_unit/wishbone_master/N2992 ;
    wire syn182169;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/C354/C3/C1 ;
    wire \bridge/pci_mux_mas_load_in ;
    wire syn20493;
    wire syn181290;
    wire syn19407;
    wire \bridge/pci_target_unit/pcit_sm_bc0_out ;
    wire syn19933;
    wire syn179287;
    wire \bridge/pci_target_unit/pcit_if_disconect_wo_data_out ;
    wire \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg ;
    wire syn181303;
    wire \bridge/output_backup/mas_ad_en_out ;
    wire \bridge/pci_mux_par_en_in ;
    wire \bridge/out_bckp_par_en_out ;
    wire syn181316;
    wire syn181329;
    wire ACK_I;
    wire syn17090;
    wire \bridge/pci_target_unit/fifos/pcir_write_performed ;
    wire syn16939;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/frame_en_slow ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/frame_en_keep ;
    wire \bridge/pci_mux_frame_en_in ;
    wire \bridge/out_bckp_frame_en_out ;
    wire \bridge/pci_target_unit/wishbone_master/C104/N6 ;
    wire syn17006;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/last_load ;
    wire syn18919;
    wire syn178584;
    wire \bridge/wishbone_slave_unit/pcim_if_last_out ;
    wire N12082;
    wire CRT_CLK_BUFGPed;
    wire \CRT/ssvga_fifo/rd_ssvga_en ;
    wire N12065;
    wire \CRT/ssvga_wbm_if/frame_read ;
    wire \CRT/ssvga_wbm_if/N1718 ;
    wire \CRT/ssvga_wbm_if/N1717 ;
    wire syn21738;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/timeout ;
    wire N12594;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/cell8 ;
    wire syn23093;
    wire syn23094;
    wire \CRT/ssvga_wbm_if/N1720 ;
    wire \CRT/ssvga_wbm_if/N1719 ;
    wire \CRT/ssvga_wbm_if/N1722 ;
    wire \CRT/ssvga_wbm_if/N1721 ;
    wire \CRT/ssvga_wbm_if/N1724 ;
    wire \CRT/ssvga_wbm_if/N1723 ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ;
    wire syn60043;
    wire syn60044;
    wire syn60045;
    wire syn177391;
    wire syn177380;
    wire syn177381;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect70 ;
    wire syn182488;
    wire syn18984;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty ;
    wire \CRT/ssvga_fifo/N739 ;
    wire \CRT/ssvga_fifo/N738 ;
    wire \CRT/ssvga_fifo/N741 ;
    wire \CRT/ssvga_fifo/N740 ;
    wire \CRT/ssvga_fifo/N743 ;
    wire \CRT/ssvga_fifo/N742 ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/C332/C3/C1 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ;
    wire \CRT/ssvga_fifo/N745 ;
    wire \CRT/ssvga_fifo/N744 ;
    wire syn181347;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out ;
    wire \CRT/ssvga_fifo/N747 ;
    wire \CRT/ssvga_fifo/N746 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/C310/C3/C1 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ;
    wire syn18908;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C14/N24 ;
    wire syn181285;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wclock_nempty_detect ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C14/N18 ;
    wire syn181298;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C14/N12 ;
    wire syn181311;
    wire \bridge/pci_target_unit/wishbone_master/C983 ;
    wire syn17011;
    wire syn17020;
    wire syn22790;
    wire syn182097;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C14/N6 ;
    wire syn181324;
    wire syn22805;
    wire syn182107;
    wire syn19710;
    wire syn182109;
    wire \bridge/pci_target_unit/del_sync_comp_req_pending_out ;
    wire syn19580;
    wire syn22771;
    wire \bridge/pci_target_unit/wishbone_master/C977 ;
    wire \bridge/wishbone_slave_unit/fifos/in_count_en ;
    wire \bridge/configuration/C338/N3 ;
    wire \bridge/configuration/delete_status_bit13 ;
    wire \bridge/configuration/delete_status_bit12 ;
    wire syn17678;
    wire syn19577;
    wire \bridge/wishbone_slave_unit/del_sync_req_req_pending_out ;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/do_del_request ;
    wire syn18939;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_slow ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep ;
    wire \bridge/pci_mux_mas_ad_en_in ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty ;
    wire \CRT/ssvga_wbm_if/N1516 ;
    wire \CRT/ssvga_wbm_if/N1515 ;
    wire syn182431;
    wire syn182432;
    wire syn23263;
    wire syn182435;
    wire \bridge/wishbone_slave_unit/fifos_wbw_full_out ;
    wire syn19385;
    wire syn19397;
    wire syn178884;
    wire \bridge/pci_target_unit/fifos/pciw_write_performed ;
    wire \CRT/ssvga_wbm_if/N1518 ;
    wire \CRT/ssvga_wbm_if/N1517 ;
    wire \bridge/parity_checker/serr_generate ;
    wire N_PAR;
    wire \bridge/parity_checker/non_critical_par ;
    wire \bridge/pci_mux_serr_en_in ;
    wire \bridge/parchk_sig_serr_out ;
    wire \CRT/ssvga_wbm_if/N1520 ;
    wire \CRT/ssvga_wbm_if/N1519 ;
    wire \bridge/pci_target_unit/pci_target_sm/state_backoff_reg ;
    wire \bridge/pci_target_unit/pci_target_sm/N64 ;
    wire \bridge/pci_target_unit/pci_target_sm/state_transfere_reg ;
    wire syn18930;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cbe_en_slow ;
    wire \bridge/pci_mux_cbe_en_in ;
    wire \bridge/out_bckp_cbe_en_out ;
    wire \bridge/configuration/delete_status_bit15 ;
    wire \bridge/configuration/delete_status_bit14 ;
    wire \CRT/ssvga_wbm_if/N1522 ;
    wire \CRT/ssvga_wbm_if/N1521 ;
    wire \CRT/ssvga_wbm_if/N1524 ;
    wire \CRT/ssvga_wbm_if/N1523 ;
    wire syn17018;
    wire \bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en ;
    wire \bridge/pci_target_unit/pcit_if_pcir_fifo_data_err_out ;
    wire syn24524;
    wire \bridge/pci_target_unit/pci_target_sm/S_89/cell0 ;
    wire syn19088;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect80 ;
    wire syn182406;
    wire \bridge/wishbone_slave_unit/fifos/out_count_en ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty ;
    wire \CRT/ssvga_wbm_if/N1526 ;
    wire \CRT/ssvga_wbm_if/N1525 ;
    wire N12436;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3384 ;
    wire syn181803;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3385 ;
    wire syn181810;
    wire \CRT/ssvga_wbm_if/N1528 ;
    wire \CRT/ssvga_wbm_if/N1527 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3386 ;
    wire syn181815;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3387 ;
    wire syn181820;
    wire \CRT/ssvga_wbm_if/N1530 ;
    wire \CRT/ssvga_wbm_if/N1529 ;
    wire N12542;
    wire \bridge/pci_target_unit/del_sync/comp_done_reg_main ;
    wire \bridge/pci_target_unit/del_sync/comp_done_reg_clr ;
    wire \bridge/pciu_pci_drcomp_pending_out ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3388 ;
    wire syn181825;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3389 ;
    wire syn181830;
    wire \CRT/ssvga_wbm_if/N1531 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3390 ;
    wire syn181835;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3391 ;
    wire syn181840;
    wire \bridge/wishbone_slave_unit/wishbone_slave/mrl_en ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/pref_en ;
    wire N12541;
    wire \bridge/pci_target_unit/del_sync/sync_req_comp_pending ;
    wire \bridge/pci_target_unit/pci_target_if/S_198/cell0 ;
    wire N12380;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C707 ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C749 ;
    wire syn16935;
    wire syn181420;
    wire \bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending ;
    wire syn22126;
    wire syn19590;
    wire syn182037;
    wire syn182038;
    wire \bridge/pci_target_unit/del_sync_comp_flush_out ;
    wire \bridge/pci_target_unit/fifos_pciw_transaction_ready_out ;
    wire \bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_done ;
    wire syn182662;
    wire syn182663;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_95/cell0 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_full ;
    wire N_LED;
    wire syn48756;
    wire syn179587;
    wire \CRT/ssvga_crtc/N400 ;
    wire syn20304;
    wire \CRT/ssvga_fifo/sync_ssvga_en ;
    wire \bridge/conf_wb_mem_io1_out ;
    wire syn176975;
    wire \CRT/ssvga_crtc/N401 ;
    wire \CRT/ssvga_crtc/N403 ;
    wire \CRT/ssvga_crtc/N402 ;
    wire \CRT/ssvga_crtc/N405 ;
    wire \CRT/ssvga_crtc/N404 ;
    wire \CRT/ssvga_crtc/N407 ;
    wire \CRT/ssvga_crtc/N406 ;
    wire \CRT/ssvga_crtc/N409 ;
    wire \CRT/ssvga_crtc/N408 ;
    wire syn17093;
    wire syn179261;
    wire \bridge/pci_target_unit/pci_target_sm/ctrl_en_w ;
    wire \bridge/pciu_pciif_devsel_en_out ;
    wire \bridge/out_bckp_trdy_en_out ;
    wire \CRT/ssvga_wbm_if/N1726 ;
    wire \CRT/ssvga_wbm_if/N1725 ;
    wire \CRT/ssvga_wbm_if/N1736 ;
    wire \CRT/ssvga_wbm_if/N1735 ;
    wire \CRT/ssvga_wbm_if/N1728 ;
    wire \CRT/ssvga_wbm_if/N1727 ;
    wire \bridge/parity_checker/par_cbe_out ;
    wire \bridge/parity_checker/cbe_par_calc/syn118 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr ;
    wire \bridge/parity_checker/cbe_par_reg ;
    wire \CRT/ssvga_wbm_if/N1746 ;
    wire \CRT/ssvga_wbm_if/N1745 ;
    wire \CRT/ssvga_wbm_if/N1738 ;
    wire \CRT/ssvga_wbm_if/N1737 ;
    wire \CRT/ssvga_wbm_if/N1730 ;
    wire \CRT/ssvga_wbm_if/N1729 ;
    wire \CRT/ssvga_wbm_if/N1740 ;
    wire \CRT/ssvga_wbm_if/N1739 ;
    wire \CRT/ssvga_wbm_if/N1732 ;
    wire \CRT/ssvga_wbm_if/N1731 ;
    wire \CRT/ssvga_wbm_if/N1742 ;
    wire \CRT/ssvga_wbm_if/N1741 ;
    wire \CRT/ssvga_wbm_if/N1734 ;
    wire \CRT/ssvga_wbm_if/N1733 ;
    wire \CRT/ssvga_wbm_if/N1744 ;
    wire \CRT/ssvga_wbm_if/N1743 ;
    wire syn17017;
    wire syn60038;
    wire \bridge/wishbone_slave_unit/del_sync_comp_req_pending_out ;
    wire syn19075;
    wire N12426;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/S_176/cell0 ;
    wire syn181630;
    wire \bridge/pci_target_unit/del_sync/req_comp_pending_sample ;
    wire N_PERR;
    wire \bridge/parity_checker/check_perr ;
    wire \bridge/parity_checker/perr_sampled ;
    wire \bridge/configuration/delete_status_bit11 ;
    wire \bridge/configuration/delete_status_bit8 ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0 ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wclock_nempty_detect90 ;
    wire syn182601;
    wire syn182602;
    wire syn182526;
    wire syn182527;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect85 ;
    wire syn182473;
    wire syn182474;
    wire syn182475;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect ;
    wire syn182394;
    wire syn182395;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect ;
    wire syn182679;
    wire syn182680;
    wire syn182682;
    wire \bridge/pci_target_unit/fifos_pciw_two_left_out ;
    wire N12162;
    wire syn16986;
    wire syn16982;
    wire syn16988;
    wire \CRT/crtc_vblank ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty ;
    wire syn182627;
    wire syn182628;
    wire syn182630;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty ;
    wire \bridge/pci_mux_frame_load_in ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame ;
    wire N12587;
    wire \bridge/pci_mux_frame_in ;
    wire \bridge/pci_target_unit/fifos/out_count_en ;
    wire syn19420;
    wire syn182538;
    wire \bridge/pci_target_unit/fifos/portA_enable ;
    wire \CRT/crtc_hblank ;
    wire \CRT/go ;
    wire \CRT/drive_blank_reg ;
    wire \bridge/out_bckp_trdy_out ;
    wire \bridge/pci_target_unit/pcit_if_read_completed_out ;
    wire syn19366;
    wire \bridge/pci_target_unit/del_sync/N1235 ;
    wire \bridge/wishbone_slave_unit/del_sync/N140 ;
    wire N12237;
    wire \bridge/wishbone_slave_unit/pcim_sm_mabort_out ;
    wire \bridge/pci_target_unit/del_sync/N1238 ;
    wire \bridge/pci_target_unit/del_sync/N1237 ;
    wire \bridge/wishbone_slave_unit/del_sync/N143 ;
    wire \bridge/wishbone_slave_unit/del_sync/N142 ;
    wire syn181426;
    wire \bridge/pci_target_unit/del_sync/N1240 ;
    wire \bridge/pci_target_unit/del_sync/N1239 ;
    wire \bridge/wishbone_slave_unit/del_sync/N145 ;
    wire \bridge/wishbone_slave_unit/del_sync/N144 ;
    wire \CRT/ssvga_wbm_if/S_41/cell0 ;
    wire syn177324;
    wire syn22076;
    wire syn21870;
    wire \bridge/pci_target_unit/del_sync/N1242 ;
    wire \bridge/pci_target_unit/del_sync/N1241 ;
    wire \bridge/wishbone_slave_unit/del_sync/N147 ;
    wire \bridge/wishbone_slave_unit/del_sync/N146 ;
    wire \bridge/pci_target_unit/del_sync/N1244 ;
    wire \bridge/pci_target_unit/del_sync/N1243 ;
    wire \bridge/wishbone_slave_unit/del_sync/N149 ;
    wire \bridge/wishbone_slave_unit/del_sync/N148 ;
    wire syn180240;
    wire syn180247;
    wire syn180248;
    wire syn20807;
    wire syn20817;
    wire syn180261;
    wire \bridge/output_backup/C3/N66 ;
    wire syn180270;
    wire syn20835;
    wire syn20841;
    wire \bridge/output_backup/C3/N72 ;
    wire syn180706;
    wire syn180707;
    wire syn180719;
    wire syn181260;
    wire syn21197;
    wire syn180720;
    wire \bridge/output_backup/C3/N126 ;
    wire syn17101;
    wire syn20872;
    wire syn20874;
    wire syn20882;
    wire syn180336;
    wire syn180337;
    wire \bridge/output_backup/C3/N78 ;
    wire syn180752;
    wire syn180753;
    wire syn180765;
    wire syn21235;
    wire syn180766;
    wire \bridge/output_backup/C3/N132 ;
    wire syn17120;
    wire syn20909;
    wire syn180385;
    wire syn20913;
    wire syn20922;
    wire syn180387;
    wire syn180388;
    wire \bridge/output_backup/C3/N84 ;
    wire syn21585;
    wire syn181217;
    wire syn181218;
    wire syn21601;
    wire syn181220;
    wire \bridge/output_backup/C3/N186 ;
    wire syn180806;
    wire syn21259;
    wire syn21274;
    wire syn180811;
    wire \bridge/output_backup/C3/N138 ;
    wire syn20947;
    wire syn180439;
    wire syn180440;
    wire syn20963;
    wire syn180442;
    wire \bridge/output_backup/C3/N90 ;
    wire syn21625;
    wire syn181272;
    wire syn181273;
    wire syn21641;
    wire syn181275;
    wire \bridge/output_backup/C3/N192 ;
    wire syn16916;
    wire syn21298;
    wire syn180855;
    wire syn21307;
    wire syn21313;
    wire \bridge/output_backup/C3/N144 ;
    wire syn20987;
    wire syn180489;
    wire syn180490;
    wire syn21003;
    wire syn180492;
    wire \bridge/output_backup/C3/N96 ;
    wire syn180899;
    wire syn21346;
    wire syn21354;
    wire syn180906;
    wire syn180907;
    wire \bridge/output_backup/C3/N150 ;
    wire syn180528;
    wire syn180529;
    wire syn180535;
    wire syn21035;
    wire syn21041;
    wire \bridge/output_backup/C3/N102 ;
    wire syn180951;
    wire syn21385;
    wire syn21396;
    wire syn180960;
    wire syn180961;
    wire \bridge/output_backup/C3/N156 ;
    wire syn180569;
    wire syn180570;
    wire syn180582;
    wire syn21080;
    wire syn180583;
    wire \bridge/output_backup/C3/N108 ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ;
    wire syn180971;
    wire syn21430;
    wire syn21436;
    wire \bridge/output_backup/C3/N162 ;
    wire syn180623;
    wire syn21104;
    wire syn21119;
    wire syn180628;
    wire \bridge/output_backup/C3/N114 ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w_frm ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy ;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_trdy_critical/syn71 ;
    wire N12472;
    wire syn180373;
    wire syn180374;
    wire syn21462;
    wire syn21479;
    wire syn181062;
    wire \bridge/output_backup/C3/N168 ;
    wire syn21143;
    wire syn180672;
    wire syn21152;
    wire syn21158;
    wire \bridge/output_backup/C3/N120 ;
    wire \bridge/pci_mux_tar_ad_en_in ;
    wire \bridge/pci_target_unit/pci_target_sm/ad_en_w ;
    wire N12338;
    wire syn181107;
    wire syn21511;
    wire syn21520;
    wire syn181113;
    wire syn181114;
    wire \bridge/output_backup/C3/N174 ;
    wire syn23454;
    wire syn181158;
    wire syn21552;
    wire syn21560;
    wire syn181165;
    wire syn181166;
    wire \bridge/output_backup/C3/N180 ;
    wire syn181508;
    wire syn181509;
    wire syn181510;
    wire syn181511;
    wire syn181520;
    wire syn181521;
    wire syn181522;
    wire syn181523;
    wire \bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit ;
    wire syn178711;
    wire syn178714;
    wire syn181624;
    wire syn19085;
    wire \bridge/parity_checker/syn415 ;
    wire \bridge/parity_checker/perr_generate ;
    wire N12031;
    wire \bridge/out_bckp_perr_out ;
    wire syn177213;
    wire \CRT/pal_wr_en ;
    wire N12543;
    wire \bridge/pci_target_unit/del_sync/sync_comp_req_pending ;
    wire N12382;
    wire syn22093;
    wire syn22095;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending ;
    wire syn22096;
    wire N12544;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_reg ;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_clr ;
    wire N12383;
    wire syn181402;
    wire syn181403;
    wire \bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_progress ;
    wire syn178847;
    wire syn178850;
    wire syn178848;
    wire syn178849;
    wire syn178853;
    wire \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg ;
    wire \bridge/pci_target_unit/pcit_sm_rdy_out ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_control_out[2] ;
    wire \bridge/parity_checker/frame_dec2 ;
    wire \CRT/ssvga_fifo/S_45/cell0 ;
    wire \CRT/ssvga_fifo/C6/N48 ;
    wire \bridge/pci_target_unit/wishbone_master/C1183 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3392 ;
    wire syn181845;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3393 ;
    wire syn181850;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3402 ;
    wire syn181895;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3394 ;
    wire syn181855;
    wire \bridge/conf_perr_response_out ;
    wire \bridge/parity_checker/pci_perr_en_reg ;
    wire N12029;
    wire \bridge/out_bckp_serr_out ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3403 ;
    wire syn181900;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3395 ;
    wire syn181860;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3412 ;
    wire syn181945;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3404 ;
    wire syn181905;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3396 ;
    wire syn181865;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3413 ;
    wire syn181950;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3405 ;
    wire syn181910;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3397 ;
    wire syn181870;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3406 ;
    wire syn181915;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3398 ;
    wire syn181875;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3407 ;
    wire syn181920;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3399 ;
    wire syn181880;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3408 ;
    wire syn181925;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3400 ;
    wire syn181885;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3409 ;
    wire syn181930;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3401 ;
    wire syn181890;
    wire N12466;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3190 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C188 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3410 ;
    wire syn181935;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3411 ;
    wire syn181940;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3193 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3192 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3195 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3194 ;
    wire syn22189;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3197 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3196 ;
    wire syn181605;
    wire syn181606;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_bound ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3191 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3198 ;
    wire \CRT/fifo_wr_en ;
    wire syn179377;
    wire syn179378;
    wire syn179382;
    wire \CRT/ssvga_fifo/S_28/cell0 ;
    wire syn20069;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_from_fifo ;
    wire \bridge/pci_target_unit/pci_target_sm/wr_to_fifo ;
    wire N12152;
    wire syn179548;
    wire syn179572;
    wire \CRT/ssvga_crtc/N326 ;
    wire \CRT/ssvga_crtc/cell25 ;
    wire \CRT/ssvga_crtc/N327 ;
    wire \CRT/ssvga_crtc/N329 ;
    wire \CRT/ssvga_crtc/N328 ;
    wire \CRT/ssvga_crtc/N331 ;
    wire \CRT/ssvga_crtc/N330 ;
    wire \CRT/ssvga_crtc/N333 ;
    wire \CRT/ssvga_crtc/N332 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 ;
    wire syn19064;
    wire \CRT/ssvga_crtc/N335 ;
    wire \CRT/ssvga_crtc/N334 ;
    wire \CRT/ssvga_fifo/S_43/cell0 ;
    wire syn20013;
    wire \bridge/in_reg_trdy_out ;
    wire \bridge/in_reg_devsel_out ;
    wire N12092;
    wire \CRT/ssvga_fifo/N801 ;
    wire \CRT/ssvga_fifo/N800 ;
    wire \bridge/pci_target_unit/pci_target_sm/devs_w ;
    wire \bridge/pci_target_unit/pci_target_sm/devs_w_frm ;
    wire \bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy ;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_devsel_critical/syn71 ;
    wire N12474;
    wire \bridge/out_bckp_devsel_out ;
    wire \CRT/ssvga_fifo/N803 ;
    wire \CRT/ssvga_fifo/N802 ;
    wire \CRT/ssvga_fifo/N805 ;
    wire \CRT/ssvga_fifo/N804 ;
    wire \CRT/ssvga_fifo/N807 ;
    wire \CRT/ssvga_fifo/N806 ;
    wire syn17012;
    wire syn17035;
    wire syn19914;
    wire syn19918;
    wire \bridge/pci_target_unit/pci_target_sm/N59 ;
    wire \bridge/pci_target_unit/pci_target_sm/previous_frame ;
    wire syn17031;
    wire syn19380;
    wire syn178869;
    wire syn179315;
    wire syn19968;
    wire syn24519;
    wire syn179246;
    wire syn179247;
    wire syn179248;
    wire syn179249;
    wire syn179245;
    wire syn19865;
    wire syn177518;
    wire syn177519;
    wire syn177524;
    wire syn177533;
    wire syn17836;
    wire syn177532;
    wire syn177514;
    wire syn177515;
    wire \bridge/configuration/C2354 ;
    wire \bridge/configuration/C2340 ;
    wire \bridge/configuration/C2308 ;
    wire syn17813;
    wire syn177511;
    wire \bridge/configuration/C2370 ;
    wire \bridge/configuration/C2338 ;
    wire syn177470;
    wire syn50321;
    wire syn177541;
    wire syn60046;
    wire syn60047;
    wire syn60048;
    wire syn60049;
    wire \bridge/configuration/C3488 ;
    wire syn177563;
    wire syn177403;
    wire syn84030;
    wire syn177475;
    wire syn177485;
    wire syn177480;
    wire \bridge/configuration/C2356 ;
    wire syn120377;
    wire syn177517;
    wire syn177508;
    wire syn177509;
    wire syn177512;
    wire syn58393;
    wire syn177632;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/C0/C116 ;
    wire syn17811;
    wire syn17815;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/C0/C108 ;
    wire syn177501;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/C0/C112 ;
    wire \bridge/configuration/C2322 ;
    wire syn177440;
    wire syn60060;
    wire syn177450;
    wire syn177451;
    wire \bridge/configuration/icr_soft_res ;
    wire \bridge/configuration/C2302 ;
    wire \bridge/configuration/C2292 ;
    wire syn177458;
    wire syn177465;
    wire \bridge/configuration/C2368 ;
    wire \bridge/configuration/C2360 ;
    wire \bridge/configuration/C2320 ;
    wire syn17049;
    wire syn177435;
    wire syn59929;
    wire syn177446;
    wire syn178109;
    wire syn16928;
    wire syn177416;
    wire syn24326;
    wire syn177631;
    wire syn16930;
    wire syn59978;
    wire syn60030;
    wire syn177580;
    wire syn177581;
    wire syn177585;
    wire syn177586;
    wire syn16917;
    wire syn17051;
    wire syn17875;
    wire syn48759;
    wire syn177570;
    wire syn177571;
    wire \bridge/configuration/C2304 ;
    wire syn177568;
    wire syn177542;
    wire syn177572;
    wire syn177573;
    wire syn177574;
    wire syn17856;
    wire syn177569;
    wire \bridge/configuration/C2334 ;
    wire syn177548;
    wire syn177393;
    wire syn177616;
    wire syn177620;
    wire syn177624;
    wire syn177625;
    wire syn17052;
    wire syn17912;
    wire syn17895;
    wire syn177611;
    wire syn177608;
    wire syn177565;
    wire \bridge/configuration/C2318 ;
    wire syn177613;
    wire syn177614;
    wire syn177617;
    wire syn17894;
    wire syn177609;
    wire syn177664;
    wire syn177665;
    wire syn177672;
    wire syn177669;
    wire syn177670;
    wire syn177656;
    wire syn177657;
    wire syn177661;
    wire syn177654;
    wire syn177655;
    wire syn177658;
    wire syn177662;
    wire syn17083;
    wire syn177629;
    wire syn50278;
    wire syn177703;
    wire syn177704;
    wire syn177705;
    wire syn17990;
    wire syn177693;
    wire syn177701;
    wire syn177710;
    wire syn177711;
    wire syn17971;
    wire syn177698;
    wire syn177699;
    wire syn177692;
    wire syn177694;
    wire syn17054;
    wire syn177743;
    wire syn177744;
    wire syn177749;
    wire syn177750;
    wire syn17115;
    wire syn177740;
    wire syn177732;
    wire syn177734;
    wire syn17055;
    wire syn177737;
    wire syn177738;
    wire syn177741;
    wire syn18010;
    wire syn177733;
    wire syn50276;
    wire syn177780;
    wire syn177781;
    wire syn177785;
    wire syn177778;
    wire syn177779;
    wire syn177782;
    wire syn177790;
    wire syn177791;
    wire syn18048;
    wire syn177822;
    wire syn177826;
    wire syn177830;
    wire syn177831;
    wire syn17057;
    wire syn18104;
    wire syn18087;
    wire syn177817;
    wire syn177814;
    wire syn177819;
    wire syn177820;
    wire syn177823;
    wire syn18086;
    wire syn177815;
    wire syn177864;
    wire syn177865;
    wire syn177870;
    wire syn17058;
    wire syn177869;
    wire syn177856;
    wire syn177857;
    wire syn177861;
    wire syn177863;
    wire syn177855;
    wire syn177858;
    wire syn177838;
    wire \bridge/configuration/config_addr[23] ;
    wire \bridge/configuration/C2296 ;
    wire syn177842;
    wire syn177897;
    wire syn177898;
    wire syn177903;
    wire syn177902;
    wire syn177889;
    wire syn177890;
    wire syn177894;
    wire syn177896;
    wire syn177888;
    wire syn177891;
    wire syn177875;
    wire \bridge/configuration/config_addr[22] ;
    wire syn17059;
    wire syn177930;
    wire syn177931;
    wire syn177936;
    wire syn177921;
    wire syn177922;
    wire syn177927;
    wire syn177923;
    wire syn177924;
    wire syn177925;
    wire syn177928;
    wire syn177935;
    wire syn17060;
    wire syn177963;
    wire syn177964;
    wire syn177969;
    wire syn177954;
    wire syn177955;
    wire syn177960;
    wire syn177956;
    wire syn177957;
    wire syn177958;
    wire syn177961;
    wire syn177968;
    wire syn17061;
    wire syn177997;
    wire syn177998;
    wire syn178003;
    wire syn17062;
    wire syn178002;
    wire syn177989;
    wire syn177990;
    wire syn177994;
    wire syn177996;
    wire syn177988;
    wire syn177991;
    wire syn177975;
    wire \bridge/configuration/config_addr[19] ;
    wire syn178030;
    wire syn178031;
    wire syn178036;
    wire syn178035;
    wire syn178022;
    wire syn178023;
    wire syn178027;
    wire syn178029;
    wire syn178021;
    wire syn178024;
    wire syn178008;
    wire \bridge/configuration/config_addr[18] ;
    wire syn17063;
    wire syn178063;
    wire syn178064;
    wire syn178069;
    wire syn178054;
    wire syn178055;
    wire syn178060;
    wire syn178056;
    wire syn178057;
    wire syn178058;
    wire syn178061;
    wire syn178068;
    wire syn17064;
    wire syn178101;
    wire syn178102;
    wire syn178107;
    wire syn17065;
    wire syn17118;
    wire syn178106;
    wire syn178092;
    wire syn178093;
    wire syn178098;
    wire syn178094;
    wire syn178095;
    wire syn178096;
    wire syn178099;
    wire syn178071;
    wire syn17772;
    wire syn178139;
    wire syn178140;
    wire syn178145;
    wire syn18431;
    wire syn178144;
    wire syn178131;
    wire syn178132;
    wire syn178136;
    wire syn178138;
    wire syn178130;
    wire syn178133;
    wire syn178117;
    wire \bridge/configuration/config_addr[15] ;
    wire syn17066;
    wire syn17067;
    wire syn178174;
    wire syn178175;
    wire syn178180;
    wire syn18468;
    wire syn178179;
    wire syn178166;
    wire syn178167;
    wire syn178171;
    wire syn178173;
    wire syn178165;
    wire syn178168;
    wire syn178152;
    wire \bridge/configuration/config_addr[14] ;
    wire syn17068;
    wire syn18511;
    wire syn178216;
    wire syn178213;
    wire syn178214;
    wire syn178205;
    wire syn178206;
    wire syn178207;
    wire syn178208;
    wire syn178200;
    wire syn178201;
    wire syn178202;
    wire syn18491;
    wire syn178204;
    wire \bridge/configuration/config_addr[13] ;
    wire syn178245;
    wire syn178246;
    wire syn178251;
    wire syn18543;
    wire syn178250;
    wire syn178236;
    wire syn178237;
    wire syn178242;
    wire syn178238;
    wire syn178239;
    wire syn178240;
    wire syn178243;
    wire syn18567;
    wire syn178265;
    wire syn178266;
    wire syn178268;
    wire syn17072;
    wire syn17071;
    wire syn17075;
    wire \bridge/configuration/config_addr[11] ;
    wire syn17073;
    wire syn17076;
    wire syn24466;
    wire syn178293;
    wire syn178294;
    wire syn178295;
    wire syn16984;
    wire syn18585;
    wire syn178292;
    wire syn17077;
    wire syn17081;
    wire syn16936;
    wire \bridge/configuration/config_addr[10] ;
    wire syn17078;
    wire syn17079;
    wire syn24468;
    wire syn178312;
    wire syn178313;
    wire syn178314;
    wire syn17119;
    wire syn178311;
    wire syn178309;
    wire syn17074;
    wire syn17080;
    wire syn24470;
    wire syn178340;
    wire syn178341;
    wire syn178342;
    wire syn178334;
    wire syn178338;
    wire syn178335;
    wire syn18636;
    wire syn17084;
    wire syn178337;
    wire \bridge/conf_pci_err_pending_out ;
    wire \bridge/conf_serr_enable_out ;
    wire syn18632;
    wire syn18633;
    wire \bridge/configuration/config_addr[8] ;
    wire syn18659;
    wire syn178356;
    wire syn178357;
    wire syn178358;
    wire syn18655;
    wire syn18658;
    wire syn24472;
    wire syn178375;
    wire syn178376;
    wire syn178377;
    wire syn18681;
    wire syn178373;
    wire syn178372;
    wire syn18670;
    wire syn24474;
    wire syn178393;
    wire syn178394;
    wire syn178395;
    wire \bridge/configuration/config_addr[5] ;
    wire syn178392;
    wire syn178390;
    wire syn18717;
    wire syn178409;
    wire syn178410;
    wire syn178411;
    wire syn18713;
    wire syn18716;
    wire syn24476;
    wire syn178435;
    wire syn178436;
    wire syn178437;
    wire syn178432;
    wire syn178433;
    wire syn18725;
    wire \bridge/configuration/serr_int_en ;
    wire syn18765;
    wire syn178470;
    wire syn18756;
    wire syn178465;
    wire syn178459;
    wire syn178460;
    wire syn178462;
    wire \bridge/configuration/wb_img_ctrl1[2] ;
    wire \bridge/configuration/perr_int_en ;
    wire \bridge/configuration/C2326 ;
    wire syn178449;
    wire syn18800;
    wire syn178494;
    wire syn178495;
    wire syn18784;
    wire syn178488;
    wire syn178489;
    wire syn178485;
    wire \bridge/configuration/error_int_en ;
    wire syn178486;
    wire syn178522;
    wire syn178523;
    wire syn178532;
    wire syn178528;
    wire syn178529;
    wire syn178530;
    wire \bridge/configuration/pci_error_en ;
    wire syn178517;
    wire syn178520;
    wire syn178516;
    wire syn17085;
    wire N12607;
    wire syn17008;
    wire syn18944;
    wire \bridge/wishbone_slave_unit/fifos/C6/N35 ;
    wire syn17669;
    wire syn177343;
    wire syn177406;
    wire syn177319;
    wire syn177320;
    wire syn177321;
    wire syn176894;
    wire syn176895;
    wire syn177317;
    wire syn177311;
    wire syn177315;
    wire syn18959;
    wire \bridge/wishbone_slave_unit/fifos/C6/N30 ;
    wire syn18965;
    wire syn18966;
    wire \bridge/wishbone_slave_unit/fifos/C6/N24 ;
    wire syn18972;
    wire syn18973;
    wire \bridge/wishbone_slave_unit/fifos/C6/N18 ;
    wire syn18979;
    wire syn18980;
    wire \bridge/wishbone_slave_unit/fifos/C6/N12 ;
    wire syn18985;
    wire \bridge/wishbone_slave_unit/fifos/C6/N6 ;
    wire syn17000;
    wire syn178898;
    wire syn178911;
    wire \bridge/pci_target_unit/fifos/C9/N30 ;
    wire syn178919;
    wire \bridge/pci_target_unit/fifos/C9/N24 ;
    wire syn178927;
    wire \bridge/pci_target_unit/fifos/C9/N18 ;
    wire syn178935;
    wire \bridge/pci_target_unit/fifos/C9/N12 ;
    wire syn178943;
    wire \bridge/pci_target_unit/fifos/C9/N6 ;
    wire syn19873;
    wire syn19881;
    wire syn19884;
    wire \bridge/conf_mem_space_enable_out ;
    wire \bridge/conf_io_space_enable_out ;
    wire \bridge/conf_pci_mem_io1_out ;
    wire \bridge/pci_target_unit/pci_target_sm/cnf_progress ;
    wire syn19963;
    wire syn17686;
    wire syn177358;
    wire \bridge/configuration/C2001 ;
    wire syn16914;
    wire syn60111;
    wire syn179659;
    wire syn20480;
    wire syn17104;
    wire syn180052;
    wire syn180053;
    wire syn180054;
    wire syn17105;
    wire syn17121;
    wire syn180051;
    wire syn17016;
    wire syn17102;
    wire \bridge/configuration/C1929 ;
    wire syn17002;
    wire syn20739;
    wire syn20740;
    wire syn20741;
    wire syn20742;
    wire syn16985;
    wire syn59991;
    wire \bridge/configuration/C1935 ;
    wire syn17003;
    wire syn17015;
    wire \bridge/configuration/C1937 ;
    wire syn17014;
    wire \bridge/configuration/C1967 ;
    wire syn17103;
    wire syn20796;
    wire syn180244;
    wire \bridge/configuration/C1941 ;
    wire syn60089;
    wire \bridge/configuration/pci_error_rty_exp_set ;
    wire \bridge/configuration/C1973 ;
    wire syn20803;
    wire syn180245;
    wire syn20934;
    wire syn48754;
    wire syn180416;
    wire syn180425;
    wire syn180417;
    wire syn180418;
    wire syn180419;
    wire syn180420;
    wire \bridge/configuration/C1989 ;
    wire \bridge/configuration/C1987 ;
    wire \bridge/configuration/C2003 ;
    wire \bridge/configuration/C1971 ;
    wire syn20953;
    wire syn16929;
    wire syn60090;
    wire syn20974;
    wire syn180466;
    wire syn180475;
    wire syn180467;
    wire syn180468;
    wire syn180469;
    wire syn180470;
    wire syn20993;
    wire syn180532;
    wire syn180534;
    wire syn16927;
    wire syn60110;
    wire syn180581;
    wire syn180580;
    wire syn16919;
    wire syn16931;
    wire syn21130;
    wire syn180657;
    wire syn180666;
    wire syn180658;
    wire syn180659;
    wire syn180660;
    wire syn180661;
    wire syn180669;
    wire syn180671;
    wire syn180718;
    wire syn180717;
    wire syn180764;
    wire syn180763;
    wire syn21285;
    wire syn180840;
    wire syn180849;
    wire syn180841;
    wire syn180842;
    wire syn180843;
    wire syn180844;
    wire syn180854;
    wire syn180852;
    wire syn21421;
    wire syn181008;
    wire syn180994;
    wire syn180995;
    wire syn181000;
    wire syn181001;
    wire syn180996;
    wire syn21407;
    wire syn180992;
    wire syn180993;
    wire \bridge/configuration/C1955 ;
    wire \bridge/configuration/C1953 ;
    wire syn17004;
    wire \bridge/configuration/C2268 ;
    wire syn181007;
    wire syn181005;
    wire syn181195;
    wire syn181196;
    wire syn181201;
    wire syn181202;
    wire syn21571;
    wire syn181193;
    wire syn181194;
    wire syn181197;
    wire syn17098;
    wire syn21589;
    wire syn181247;
    wire syn181248;
    wire syn181253;
    wire syn181258;
    wire syn181249;
    wire syn181250;
    wire syn181251;
    wire syn181252;
    wire syn21629;
    wire syn181498;
    wire syn181499;
    wire syn181512;
    wire syn181497;
    wire syn176956;
    wire syn176958;
    wire syn181495;
    wire syn181500;
    wire syn181501;
    wire syn181502;
    wire syn181503;
    wire syn176967;
    wire syn176960;
    wire syn176963;
    wire syn176965;
    wire syn181504;
    wire syn181505;
    wire syn181506;
    wire syn181507;
    wire syn176969;
    wire syn176971;
    wire syn176973;
    wire syn176977;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/C0/C104 ;
    wire syn182355;
    wire \bridge/pci_target_unit/pci_target_sm/load_med_reg_w ;
    wire \bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy ;
    wire syn19415;
    wire \bridge/pci_target_unit/pcit_sm_load_medium_reg_out ;
    wire syn17010;
    wire syn178535;
    wire syn178547;
    wire syn177332;
    wire syn17053;
    wire syn18051;
    wire syn177771;
    wire syn177772;
    wire syn177773;
    wire syn17070;
    wire syn178514;
    wire syn178515;
    wire syn178518;
    wire syn17087;
    wire syn178727;
    wire syn17086;
    wire \bridge/wishbone_slave_unit/fifos/C3/N30 ;
    wire syn19081;
    wire syn178708;
    wire syn178718;
    wire syn178732;
    wire \bridge/wishbone_slave_unit/fifos/C3/N24 ;
    wire syn178737;
    wire \bridge/wishbone_slave_unit/fifos/C3/N18 ;
    wire syn178742;
    wire \bridge/wishbone_slave_unit/fifos/C3/N12 ;
    wire syn178747;
    wire \bridge/wishbone_slave_unit/fifos/C3/N6 ;
    wire syn178873;
    wire syn179034;
    wire \bridge/pci_target_unit/fifos/C10/N30 ;
    wire syn178998;
    wire syn178999;
    wire syn179042;
    wire \bridge/pci_target_unit/fifos/C10/N24 ;
    wire syn179050;
    wire \bridge/pci_target_unit/fifos/C10/N18 ;
    wire syn179058;
    wire \bridge/pci_target_unit/fifos/C10/N12 ;
    wire syn179066;
    wire \bridge/pci_target_unit/fifos/C10/N6 ;
    wire syn179294;
    wire syn17097;
    wire syn20373;
    wire syn20406;
    wire syn179711;
    wire \bridge/configuration/C285/N34 ;
    wire syn20389;
    wire syn20360;
    wire syn20371;
    wire syn179694;
    wire syn20359;
    wire syn179707;
    wire syn179708;
    wire syn179709;
    wire \bridge/configuration/C1959 ;
    wire \bridge/configuration/C1925 ;
    wire \bridge/configuration/C1951 ;
    wire syn179850;
    wire syn179851;
    wire syn179855;
    wire syn179846;
    wire syn179847;
    wire syn179848;
    wire syn179849;
    wire \bridge/configuration/wb_img_ctrl1[0] ;
    wire \bridge/configuration/int_prop_en ;
    wire syn179869;
    wire syn20490;
    wire syn20482;
    wire syn20484;
    wire \bridge/pci_mux_tar_load_in ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/load_force ;
    wire syn20523;
    wire syn179919;
    wire syn179920;
    wire syn179910;
    wire syn179911;
    wire syn179912;
    wire syn179913;
    wire syn179918;
    wire syn179949;
    wire syn179950;
    wire syn179954;
    wire syn179948;
    wire syn179951;
    wire syn179957;
    wire syn179959;
    wire syn179986;
    wire syn179987;
    wire syn179988;
    wire syn179989;
    wire syn179985;
    wire syn180000;
    wire syn180030;
    wire syn180031;
    wire syn180032;
    wire syn180033;
    wire syn17110;
    wire syn17111;
    wire syn17107;
    wire syn17109;
    wire syn180064;
    wire syn180081;
    wire syn180082;
    wire syn180083;
    wire syn180084;
    wire syn16983;
    wire \bridge/configuration/config_addr[6] ;
    wire syn17099;
    wire syn180095;
    wire syn180120;
    wire syn180121;
    wire syn180122;
    wire syn180123;
    wire syn180167;
    wire syn180138;
    wire syn180141;
    wire syn180205;
    wire syn180209;
    wire syn20770;
    wire syn20771;
    wire syn20772;
    wire syn20773;
    wire syn180198;
    wire syn180202;
    wire syn20769;
    wire syn180258;
    wire syn180283;
    wire syn180284;
    wire syn180285;
    wire syn180282;
    wire syn180281;
    wire syn20853;
    wire syn180313;
    wire syn180321;
    wire syn180314;
    wire syn180315;
    wire syn180316;
    wire syn180317;
    wire syn180322;
    wire syn180329;
    wire syn20893;
    wire syn180365;
    wire syn180366;
    wire syn180367;
    wire syn180368;
    wire syn180369;
    wire syn180381;
    wire syn20911;
    wire syn180432;
    wire syn180482;
    wire syn21014;
    wire syn180520;
    wire syn180521;
    wire syn180522;
    wire syn180523;
    wire syn180524;
    wire syn180500;
    wire syn180577;
    wire syn21053;
    wire syn180561;
    wire syn180562;
    wire syn180563;
    wire syn180564;
    wire syn180565;
    wire syn21091;
    wire syn180607;
    wire syn180616;
    wire syn180608;
    wire syn180609;
    wire syn180610;
    wire syn180611;
    wire syn180627;
    wire syn180626;
    wire syn180637;
    wire syn180714;
    wire syn21170;
    wire syn180698;
    wire syn180699;
    wire syn180700;
    wire syn180701;
    wire syn180702;
    wire syn180760;
    wire syn21208;
    wire syn180744;
    wire syn180745;
    wire syn180746;
    wire syn180747;
    wire syn180748;
    wire syn21246;
    wire syn180790;
    wire syn180799;
    wire syn180791;
    wire syn180792;
    wire syn180793;
    wire syn180794;
    wire syn180810;
    wire syn180809;
    wire syn180820;
    wire syn21325;
    wire syn180888;
    wire syn180892;
    wire syn180884;
    wire syn180885;
    wire syn180886;
    wire syn180887;
    wire syn180883;
    wire \bridge/configuration/status_bit8 ;
    wire syn21342;
    wire syn21365;
    wire syn180940;
    wire syn180944;
    wire syn180936;
    wire syn180937;
    wire syn180938;
    wire syn180939;
    wire syn17056;
    wire syn180935;
    wire syn180957;
    wire syn180958;
    wire syn181039;
    wire syn181040;
    wire syn181045;
    wire syn181046;
    wire syn21448;
    wire syn181037;
    wire syn181038;
    wire syn181041;
    wire syn181054;
    wire syn21465;
    wire syn21466;
    wire syn120365;
    wire syn181060;
    wire syn181058;
    wire \bridge/configuration/C2240 ;
    wire syn21490;
    wire syn181096;
    wire syn181100;
    wire syn181092;
    wire syn181093;
    wire syn181094;
    wire syn181095;
    wire syn181091;
    wire syn21506;
    wire syn21507;
    wire syn21531;
    wire syn181147;
    wire syn181151;
    wire syn181143;
    wire syn181144;
    wire syn181145;
    wire syn181146;
    wire syn181142;
    wire syn21548;
    wire syn181210;
    wire syn181265;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/tabort_ff_in ;
    wire syn22184;
    wire \bridge/wishbone_slave_unit/pcim_sm_first_out ;
    wire syn22083;
    wire \bridge/in_reg_stop_out ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C248 ;
    wire syn22101;
    wire \bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out ;
    wire syn22812;
    wire \bridge/pci_target_unit/del_sync/comp_rty_exp_reg ;
    wire syn23126;
    wire syn19708;
    wire syn19709;
    wire syn179112;
    wire syn179113;
    wire syn19701;
    wire syn19698;
    wire syn179111;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn137 ;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn129 ;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/ch_state_med ;
    wire syn177262;
    wire syn177263;
    wire syn177264;
    wire syn177265;
    wire syn176876;
    wire syn177260;
    wire syn177249;
    wire syn177253;
    wire syn177257;
    wire \CRT/ssvga_fifo/C6/N54 ;
    wire syn19959;
    wire syn20367;
    wire syn179679;
    wire syn20368;
    wire \bridge/configuration/config_addr[4] ;
    wire syn180029;
    wire \bridge/configuration/config_addr[7] ;
    wire syn180119;
    wire syn180162;
    wire syn17005;
    wire syn181111;
    wire syn181563;
    wire syn181562;
    wire \bridge/parity_checker/perr_en_crit_gen/syn112 ;
    wire N12033;
    wire \bridge/parity_checker/syn3156 ;
    wire \bridge/parity_checker/syn3166 ;
    wire \bridge/parity_checker/syn3083 ;
    wire \bridge/parity_checker/syn3174 ;
    wire \bridge/parity_checker/syn3096 ;
    wire \bridge/parity_checker/syn3164 ;
    wire \bridge/parity_checker/syn3155 ;
    wire syn18066;
    wire \bridge/wishbone_slave_unit/fifos/C3/N33 ;
    wire \bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy ;
    wire \bridge/pci_target_unit/pci_target_sm/read_completed_reg ;
    wire syn179021;
    wire \bridge/pci_target_unit/wishbone_master/C82/C0 ;
    wire N12510;
    wire syn179376;
    wire syn179379;
    wire \CRT/ssvga_crtc/line_end2 ;
    wire \CRT/ssvga_crtc/line_end1 ;
    wire syn16991;
    wire \bridge/configuration/wb_error_en ;
    wire syn16992;
    wire syn16934;
    wire syn179761;
    wire syn179762;
    wire \bridge/configuration/C281/N3 ;
    wire syn22225;
    wire syn22226;
    wire syn181988;
    wire syn181989;
    wire syn181990;
    wire syn181991;
    wire syn182000;
    wire syn182001;
    wire syn182002;
    wire syn182003;
    wire \bridge/pci_target_unit/wishbone_master/C723 ;
    wire syn23069;
    wire syn178588;
    wire \bridge/wishbone_slave_unit/del_sync_burst_out ;
    wire syn179535;
    wire N12151;
    wire \bridge/configuration/C1919 ;
    wire syn179775;
    wire syn179776;
    wire syn17043;
    wire syn17100;
    wire \bridge/configuration/C289/N9 ;
    wire syn181992;
    wire syn181993;
    wire syn181994;
    wire syn181995;
    wire syn181996;
    wire syn181997;
    wire syn181998;
    wire syn181999;
    wire syn182052;
    wire syn182285;
    wire syn23022;
    wire syn182403;
    wire syn182404;
    wire syn182423;
    wire syn182424;
    wire syn182484;
    wire syn182485;
    wire syn182486;
    wire syn182535;
    wire syn182536;
    wire syn182564;
    wire syn182565;
    wire syn182555;
    wire syn182556;
    wire syn182576;
    wire syn182577;
    wire syn182610;
    wire syn182611;
    wire syn182650;
    wire syn182651;
    wire \bridge/parity_checker/syn3204 ;
    wire \bridge/parity_checker/syn3214 ;
    wire \bridge/parity_checker/syn3125 ;
    wire \bridge/parity_checker/syn3210 ;
    wire \bridge/parity_checker/data_par ;
    wire \bridge/parity_checker/syn3203 ;
    wire syn19202;
    wire syn20277;
    wire syn179567;
    wire N12164;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/irdy_slow ;
    wire \bridge/pci_mux_irdy_in ;
    wire \bridge/pci_target_unit/pci_target_if/bckp_trdy_reg ;
    wire \bridge/pci_target_unit/pci_target_if/trdy_asserted_reg ;
    wire N12540;
    wire \bridge/pci_target_unit/del_sync/req_done_reg ;
    wire \bridge/configuration/C299/N74 ;
    wire \bridge/configuration/config_addr[12] ;
    wire \bridge/configuration/C299/N29 ;
    wire \bridge/configuration/config_addr[21] ;
    wire \bridge/configuration/config_addr[16] ;
    wire \bridge/configuration/config_addr[17] ;
    wire \bridge/configuration/C290/N54 ;
    wire \bridge/configuration/C290/N99 ;
    wire \bridge/configuration/config_addr[20] ;
    wire \bridge/configuration/C290/N3 ;
    wire \bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr ;
    wire \bridge/pci_target_unit/del_sync/comp_rty_exp_clr ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr ;
    wire N12313;
    wire \bridge/configuration/C299/N99 ;
    wire \bridge/configuration/config_addr[3] ;
    wire \bridge/configuration/config_addr[9] ;
    wire \bridge/configuration/C301/N3 ;
    wire \bridge/configuration/C294/N84 ;
    wire \bridge/configuration/C294/N69 ;
    wire \bridge/configuration/C294/N29 ;
    wire \bridge/pci_io_mux/ad_load_ctrl_mhigh ;
    wire \bridge/pci_io_mux/ad_load_ctrl_low ;
    wire \bridge/configuration/C291/N94 ;
    wire \bridge/configuration/C291/N59 ;
    wire \bridge/configuration/C291/N14 ;
    wire \bridge/configuration/C292/N3 ;
    wire N12330;
    wire \bridge/parity_checker/syn3190 ;
    wire \bridge/parity_checker/syn3189 ;
    wire \bridge/parity_checker/syn3172 ;
    wire \bridge/parity_checker/master_perr_report ;
    wire \bridge/parchk_par_err_detect_out ;
    wire \bridge/out_bckp_irdy_en_out ;
    wire \bridge/configuration/config_addr[2] ;
    wire \bridge/configuration/config_addr[0] ;
    wire \bridge/configuration/C296/N64 ;
    wire \bridge/configuration/C296/N89 ;
    wire \bridge/configuration/C296/N24 ;
    wire N12379;
    wire \bridge/wishbone_slave_unit/del_sync/req_done_reg ;
    wire \bridge/configuration/C346/N5 ;
    wire \bridge/configuration/delete_wb_err_cs_bit8 ;
    wire crt_hsync;
    wire \bridge/configuration/C295/N3 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/frame_load_slow ;
    wire \bridge/pci_target_unit/del_sync/sync_comp_done ;
    wire \bridge/configuration/C297/N84 ;
    wire \bridge/configuration/C297/N69 ;
    wire \bridge/configuration/C297/N29 ;
    wire \bridge/pci_io_mux/ad_load_ctrl_high ;
    wire \bridge/pci_io_mux/ad_load_ctrl_mlow ;
    wire \bridge/pci_target_unit/del_sync/sync_req_rty_exp ;
    wire \bridge/configuration/C293/N14 ;
    wire \CRT/ssvga_fifo/C6/N18 ;
    wire \CRT/ssvga_fifo/C6/N12 ;
    wire \CRT/ssvga_fifo/C6/N30 ;
    wire \CRT/ssvga_fifo/C6/N24 ;
    wire \CRT/ssvga_fifo/C6/N42 ;
    wire \CRT/ssvga_fifo/C6/N36 ;
    wire \bridge/configuration/C288/N39 ;
    wire \bridge/configuration/C283/N39 ;
    wire \bridge/configuration/C302/N19 ;
    wire \bridge/configuration/C286/N54 ;
    wire \bridge/configuration/C286/N99 ;
    wire \bridge/configuration/C286/N19 ;
    wire N12378;
    wire \bridge/wbu_mabort_rec_out ;
    wire N12381;
    wire syn120398;
    wire \CRT/ssvga_wbm_if/C1472/C18/C1/O ;
    wire syn19713;
    wire syn19562;
    wire syn178883;
    wire \bridge/pci_target_unit/pci_target_if/n_1317 ;
    wire \bridge/pci_target_unit/pci_target_if/n_1352 ;
    wire syn120402;
    wire \bridge/pci_target_unit/fifos/portB_enable ;
    wire syn120400;
    wire syn21610;
    wire \bridge/configuration/C287/N3 ;
    wire syn17023;
    wire \bridge/wishbone_slave_unit/del_sync_comp_flush_out ;
    wire \bridge/pci_target_unit/pci_target_if/N5157 ;
    wire syn120386;
    wire syn120394;
    wire syn120384;
    wire syn179789;
    wire syn120382;
    wire \bridge/pci_target_unit/pci_target_if/n_1298 ;
    wire \bridge/configuration/C284/N39 ;
    wire \bridge/pci_target_unit/pci_target_if/n_1335 ;
    wire N12539;
    wire \bridge/configuration/C285/N99 ;
    wire \bridge/configuration/C280/N3 ;
    wire \bridge/configuration/C298/N3 ;
    wire \bridge/pciu_pciif_tabort_set_out ;
    wire \bridge/configuration/C285/N79 ;
    wire syn179544;
    wire N12163;
    wire N12312;
    wire \CRT/ssvga_fifo/C6/N6 ;
    wire \bridge/parity_checker/par_out_only ;
    wire \bridge/parity_checker/par_gen/syn143 ;
    wire \bridge/pci_mux_par_in ;
    wire \bridge/parity_checker/syn3208 ;
    wire \bridge/parity_checker/syn3196 ;
    wire \bridge/parity_checker/syn3148 ;
    wire N12322;
    wire N12314;
    wire crt_vsync;
    wire \C20042/IBUFG ;
    wire \C20043/IBUFG ;
    wire GLOBAL_LOGIC0;
    wire GLOBAL_LOGIC1;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C4/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C6/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C8/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C10/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C12/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C14/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C16/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C18/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C20/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C22/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C24/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C26/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C28/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C30/C1/O ;
    wire \CRT/ssvga_fifo/C748/C4/C1/O ;
    wire \CRT/ssvga_fifo/C748/C6/C1/O ;
    wire \CRT/ssvga_fifo/C748/C8/C1/O ;
    wire \CRT/ssvga_fifo/C748/C10/C1/O ;
    wire \CRT/ssvga_wbm_if/C1472/C4/C1/O ;
    wire \CRT/ssvga_wbm_if/C1472/C6/C1/O ;
    wire \CRT/ssvga_wbm_if/C1472/C8/C1/O ;
    wire \CRT/ssvga_wbm_if/C1472/C10/C1/O ;
    wire \CRT/ssvga_wbm_if/C1472/C12/C1/O ;
    wire \CRT/ssvga_wbm_if/C1472/C14/C1/O ;
    wire \CRT/ssvga_wbm_if/C1472/C16/C1/O ;
    wire \CRT/ssvga_fifo/C749/C4/C1/O ;
    wire \CRT/ssvga_fifo/C749/C6/C1/O ;
    wire \CRT/ssvga_fifo/C749/C8/C1/O ;
    wire \bridge/pci_target_unit/del_sync/C1264/C4/C1/O ;
    wire \bridge/pci_target_unit/del_sync/C1264/C6/C1/O ;
    wire \bridge/pci_target_unit/del_sync/C1264/C8/C1/O ;
    wire \bridge/pci_target_unit/del_sync/C1264/C10/C1/O ;
    wire \bridge/pci_target_unit/del_sync/C1264/C12/C1/O ;
    wire \bridge/pci_target_unit/del_sync/C1264/C14/C1/O ;
    wire \bridge/pci_target_unit/del_sync/C1264/C16/C1/O ;
    wire \bridge/pci_target_unit/del_sync/C1264/C18/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C4/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C6/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C8/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C10/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C12/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C14/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C16/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C18/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C20/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C22/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C24/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C26/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C28/C1/O ;
    wire \CRT/ssvga_wbm_if/C1473/C30/C1/O ;
    wire \CRT/ssvga_crtc/C529/C4/C1/O ;
    wire \CRT/ssvga_crtc/C529/C6/C1/O ;
    wire \CRT/ssvga_crtc/C529/C8/C1/O ;
    wire \CRT/ssvga_crtc/C529/C10/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3410/C4/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3410/C6/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3410/C8/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C3/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C5/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C7/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C9/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C11/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C13/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C15/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C17/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C19/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C21/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C23/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C25/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C27/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C29/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C31/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3411/C4/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3110 ;
    wire \bridge/pci_target_unit/wishbone_master/N3111 ;
    wire \bridge/pci_target_unit/wishbone_master/C3411/C6/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3112 ;
    wire \bridge/pci_target_unit/wishbone_master/N3113 ;
    wire \bridge/pci_target_unit/wishbone_master/C3411/C8/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3114 ;
    wire \bridge/pci_target_unit/wishbone_master/N3115 ;
    wire \bridge/pci_target_unit/wishbone_master/N3116 ;
    wire \bridge/pci_target_unit/wishbone_master/N3117 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C4/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C6/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C8/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C4/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C6/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C8/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C10/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C12/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C14/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C16/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C18/C1/O ;
    wire \CRT/ssvga_crtc/C530/C4/C1/O ;
    wire \CRT/ssvga_crtc/C530/C6/C1/O ;
    wire \CRT/ssvga_crtc/C530/C8/C1/O ;
    wire \CRT/ssvga_crtc/C530/C10/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C4/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C6/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C8/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C10/C1/O ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/n_850 ;
    wire GLOBAL_LOGIC0_0;
    wire GLOBAL_LOGIC0_1;
    wire GLOBAL_LOGIC0_2;
    wire GLOBAL_LOGIC0_3;
    wire GLOBAL_LOGIC0_4;
    wire GLOBAL_LOGIC0_5;
    wire GLOBAL_LOGIC0_6;
    wire GLOBAL_LOGIC0_7;
    wire GLOBAL_LOGIC0_8;
    wire GLOBAL_LOGIC0_9;
    wire GLOBAL_LOGIC0_10;
    wire GLOBAL_LOGIC0_11;
    wire \bridge/configuration/delete_pci_err_cs_bit10/SRNOT ;
    wire \bridge/configuration/delete_pci_err_cs_bit10/GROM ;
    wire \bridge/configuration/C387/N3 ;
    wire \bridge/configuration/delete_pci_err_cs_bit10/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/delete_pci_err_cs_bit10/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[0]/SRNOT ;
    wire \bridge/out_bckp_ad_out[0]/GROM ;
    wire \bridge/out_bckp_ad_out[0]/FROM ;
    wire \bridge/out_bckp_ad_out[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[1]/SRNOT ;
    wire \bridge/out_bckp_ad_out[1]/GROM ;
    wire \bridge/out_bckp_ad_out[1]/FROM ;
    wire \bridge/out_bckp_ad_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[3]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[3]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[2]/SRNOT ;
    wire \bridge/out_bckp_ad_out[2]/GROM ;
    wire \bridge/out_bckp_ad_out[2]/FROM ;
    wire \bridge/out_bckp_ad_out[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[1]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C107/N5 ;
    wire \bridge/pci_target_unit/wishbone_master/C107/N10 ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[3]/SRNOT ;
    wire \bridge/out_bckp_ad_out[3]/GROM ;
    wire \bridge/out_bckp_ad_out[3]/FROM ;
    wire \bridge/out_bckp_ad_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_burst_out/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_burst_out ;
    wire \bridge/pci_target_unit/del_sync_burst_out/FROM ;
    wire \bridge/pci_target_unit/del_sync_burst_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[5]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[5]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[5]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[4]/SRNOT ;
    wire \bridge/out_bckp_ad_out[4]/GROM ;
    wire \bridge/out_bckp_ad_out[4]/FROM ;
    wire \bridge/out_bckp_ad_out[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[3]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C107/N15 ;
    wire \bridge/pci_target_unit/wishbone_master/C107/N20 ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[5]/SRNOT ;
    wire \bridge/out_bckp_ad_out[5]/GROM ;
    wire \bridge/out_bckp_ad_out[5]/FROM ;
    wire \bridge/out_bckp_ad_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[7]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[7]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[7]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[6]/SRNOT ;
    wire \bridge/out_bckp_ad_out[6]/GROM ;
    wire \bridge/out_bckp_ad_out[6]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[5]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C107/N25 ;
    wire \bridge/pci_target_unit/wishbone_master/C107/N30 ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \ADR_O[10]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N66 ;
    wire \ADR_O[10]/FROM ;
    wire \ADR_O[10]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[7]/SRNOT ;
    wire \bridge/out_bckp_ad_out[7]/GROM ;
    wire \bridge/out_bckp_ad_out[7]/FROM ;
    wire \bridge/out_bckp_ad_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[8]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[8]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[8]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[8]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[11]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N72 ;
    wire \bridge/pciu_err_addr_out[11]/FROM ;
    wire \bridge/pciu_err_addr_out[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[8]/SRNOT ;
    wire \bridge/out_bckp_ad_out[8]/GROM ;
    wire \bridge/out_bckp_ad_out[8]/FROM ;
    wire \bridge/out_bckp_ad_out[8]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[7]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C107/N35 ;
    wire \bridge/pci_target_unit/wishbone_master/C107/N40 ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/rty_counter[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[9]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[9]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[9]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[20]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N126 ;
    wire \bridge/pciu_err_addr_out[20]/FROM ;
    wire \bridge/pciu_err_addr_out[20]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[12]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N78 ;
    wire \bridge/pciu_err_addr_out[12]/FROM ;
    wire \bridge/pciu_err_addr_out[12]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[9]/SRNOT ;
    wire \bridge/out_bckp_ad_out[9]/GROM ;
    wire \bridge/out_bckp_ad_out[9]/FROM ;
    wire \bridge/out_bckp_ad_out[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[21]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N132 ;
    wire \bridge/pciu_err_addr_out[21]/FROM ;
    wire \bridge/pciu_err_addr_out[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[13]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N84 ;
    wire \bridge/pciu_err_addr_out[13]/FROM ;
    wire \bridge/pciu_err_addr_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[30]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N186 ;
    wire \bridge/pciu_err_addr_out[30]/FROM ;
    wire \bridge/pciu_err_addr_out[30]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[22]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N138 ;
    wire \bridge/pciu_err_addr_out[22]/FROM ;
    wire \bridge/pciu_err_addr_out[22]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[14]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N90 ;
    wire \bridge/pciu_err_addr_out[14]/FROM ;
    wire \bridge/pciu_err_addr_out[14]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[31]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N192 ;
    wire \bridge/pciu_err_addr_out[31]/FROM ;
    wire \bridge/pciu_err_addr_out[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[23]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N144 ;
    wire \bridge/pciu_err_addr_out[23]/FROM ;
    wire \bridge/pciu_err_addr_out[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[15]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N96 ;
    wire \bridge/pciu_err_addr_out[15]/FROM ;
    wire \bridge/pciu_err_addr_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[24]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N150 ;
    wire \bridge/pciu_err_addr_out[24]/FROM ;
    wire \bridge/pciu_err_addr_out[24]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[16]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N102 ;
    wire \bridge/pciu_err_addr_out[16]/FROM ;
    wire \bridge/pciu_err_addr_out[16]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[25]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N156 ;
    wire \bridge/pciu_err_addr_out[25]/FROM ;
    wire \bridge/pciu_err_addr_out[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[17]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N108 ;
    wire \bridge/pciu_err_addr_out[17]/FROM ;
    wire \bridge/pciu_err_addr_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[26]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N162 ;
    wire \bridge/pciu_err_addr_out[26]/FROM ;
    wire \bridge/pciu_err_addr_out[26]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[18]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N114 ;
    wire \bridge/pciu_err_addr_out[18]/FROM ;
    wire \bridge/pciu_err_addr_out[18]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N5 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_stop_out/SRNOT ;
    wire \bridge/out_bckp_stop_out/GROM ;
    wire \bridge/out_bckp_stop_out/FROM ;
    wire \bridge/out_bckp_stop_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[27]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N168 ;
    wire \bridge/pciu_err_addr_out[27]/FROM ;
    wire \bridge/pciu_err_addr_out[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[19]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N120 ;
    wire \bridge/pciu_err_addr_out[19]/FROM ;
    wire \bridge/pciu_err_addr_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N10 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N17 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[28]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N174 ;
    wire \bridge/pciu_err_addr_out[28]/FROM ;
    wire \bridge/pciu_err_addr_out[28]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_full ;
    wire \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[29]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N180 ;
    wire \bridge/pciu_err_addr_out[29]/FROM ;
    wire \bridge/pciu_err_addr_out[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N6 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N12 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[1]/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N18 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N24 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[3]/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N30 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N36 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[4]/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_raddr_0[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N42 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N48 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_rdy_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/rdy_out358 ;
    wire \bridge/wishbone_slave_unit/pcim_if_rdy_out/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_rdy_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/wr_progress/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/read_request ;
    wire \bridge/pci_target_unit/pci_target_sm/write_progress ;
    wire \bridge/pci_target_unit/pci_target_sm/wr_progress/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/wr_progress/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFX/SET ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N361 ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N362 ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N345 ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N346 ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N272 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N273 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N327 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N328 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N363 ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N347 ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[4]/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N274 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N329 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N275 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[0]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[0]/GROM ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C3/N5 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/N1961 ;
    wire \bridge/pci_target_unit/fifos/N1962 ;
    wire \bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_conf_offset_out[8]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/C19/N5 ;
    wire \bridge/pciu_conf_offset_out[8]/FROM ;
    wire \bridge/pciu_conf_offset_out[8]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_conf_offset_out[8]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[11]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[11]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[11]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[21]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[21]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[21]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[13]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[13]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[13]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[31]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[31]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[31]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[23]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[23]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[23]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[15]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[15]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[15]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[25]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[25]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[25]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[17]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[17]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[17]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_almost_full_in ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_full ;
    wire \bridge/pci_target_unit/fifos_pcir_full_out/FFY/RST ;
    wire \bridge/pci_target_unit/fifos_pcir_full_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos_pcir_full_out/FFX/RST ;
    wire \bridge/pci_target_unit/fifos_pcir_full_out/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[27]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[27]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[27]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[19]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[19]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[19]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N192 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N186 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[11]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N55 ;
    wire \bridge/pci_target_unit/del_sync/C1265/N60 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[29]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[29]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[29]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_addr_out[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N55 ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N60 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N180 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N174 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[13]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N65 ;
    wire \bridge/pci_target_unit/del_sync/C1265/N70 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/same_read_reg/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/same_read_reg/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/same_read_reg/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/same_read_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/same_read_reg/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N65 ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N70 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N168 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N162 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[15]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N75 ;
    wire \bridge/pci_target_unit/del_sync/C1265/N80 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N75 ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N80 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/SRNOT ;
    wire \CRT/ssvga_wbs_if/N40 ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N156 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N150 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[1]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N85 ;
    wire \bridge/pci_target_unit/del_sync/C1265/N10 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N85 ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N10 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N144 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N138 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[0]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N6 ;
    wire \bridge/pciu_err_addr_out[0]/FROM ;
    wire \bridge/pciu_err_addr_out[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/in_reg_idsel_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/wbs_sm_lock_in ;
    wire \bridge/in_reg_idsel_out/FROM ;
    wire \bridge/in_reg_idsel_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/in_reg_idsel_out/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_addr_out[1]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N12 ;
    wire \bridge/pciu_err_addr_out[1]/FROM ;
    wire \bridge/pciu_err_addr_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \ADR_O[2]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N18 ;
    wire \ADR_O[2]/FROM ;
    wire \ADR_O[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_cs_bit31_24[30]/SRNOT ;
    wire \bridge/configuration/pci_err_cs_bit31_24[30]/GROM ;
    wire \bridge/configuration/pci_err_cs_bit31_24[30]/FROM ;
    wire \bridge/configuration/pci_err_cs_bit31_24[30]/FFY/ASYNC_FF_GSR_OR ;
    wire \ADR_O[3]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N24 ;
    wire \ADR_O[3]/FROM ;
    wire \ADR_O[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_cs_bit31_24[31]/SRNOT ;
    wire N12518;
    wire \bridge/configuration/pci_err_cs_bit31_24[31]/FROM ;
    wire \bridge/configuration/pci_err_cs_bit31_24[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \ADR_O[4]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N30 ;
    wire \ADR_O[4]/FROM ;
    wire \ADR_O[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \ADR_O[5]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N36 ;
    wire \ADR_O[5]/FROM ;
    wire \ADR_O[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \ADR_O[6]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N42 ;
    wire \ADR_O[6]/FROM ;
    wire \ADR_O[6]/FFY/ASYNC_FF_GSR_OR ;
    wire \ADR_O[7]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N48 ;
    wire \ADR_O[7]/FROM ;
    wire \ADR_O[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \ADR_O[8]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N54 ;
    wire \ADR_O[8]/FROM ;
    wire \ADR_O[8]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_cs_bit31_24[29]/SRNOT ;
    wire \bridge/configuration/pci_err_cs_bit31_24[29]/GROM ;
    wire \bridge/configuration/pci_err_cs_bit31_24[29]/FROM ;
    wire \bridge/configuration/pci_err_cs_bit31_24[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_cs_bit31_24[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \ADR_O[9]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3415/N60 ;
    wire \ADR_O[9]/FROM ;
    wire \ADR_O[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[3]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N322 ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N323 ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[4]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N324 ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[4]/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_cbe_out[0]/SRNOT ;
    wire \bridge/out_bckp_cbe_out[0]/GROM ;
    wire \bridge/out_bckp_cbe_out[0]/FROM ;
    wire \bridge/out_bckp_cbe_out[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_cbe_out[1]/SRNOT ;
    wire \bridge/out_bckp_cbe_out[1]/GROM ;
    wire \bridge/out_bckp_cbe_out[1]/FROM ;
    wire \bridge/out_bckp_cbe_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_par_en_out/SRNOT ;
    wire \bridge/out_bckp_par_en_out/GROM ;
    wire \bridge/out_bckp_par_en_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_cbe_out[2]/SRNOT ;
    wire \bridge/out_bckp_cbe_out[2]/GROM ;
    wire \bridge/out_bckp_cbe_out[2]/FROM ;
    wire \bridge/out_bckp_cbe_out[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_cbe_out[3]/SRNOT ;
    wire \bridge/out_bckp_cbe_out[3]/GROM ;
    wire \bridge/out_bckp_cbe_out[3]/FROM ;
    wire \bridge/out_bckp_cbe_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_write_performed/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pcir_write_performed/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_write_performed/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_write_performed/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_frame_en_out/SRNOT ;
    wire \bridge/out_bckp_frame_en_out/GROM ;
    wire \bridge/out_bckp_frame_en_out/FROM ;
    wire \bridge/out_bckp_frame_en_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C103/N5 ;
    wire \bridge/pci_target_unit/wishbone_master/C103/N10 ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_last_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_next_last_out ;
    wire \bridge/wishbone_slave_unit/pcim_if_last_out/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[1]/SRNOT ;
    wire \CRT/ssvga_fifo/C2/N50 ;
    wire \CRT/ssvga_fifo/C2/N45 ;
    wire \CRT/ssvga_fifo/rd_ptr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N6 ;
    wire \CRT/ssvga_wbm_if/C1475/N12 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/timeout/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/last_transfered265 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/timeout509 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/timeout/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/timeout/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_bc_out[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C26/N6 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C26/N12 ;
    wire \bridge/wishbone_slave_unit/pcim_if_bc_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_bc_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[3]/SRNOT ;
    wire \CRT/ssvga_fifo/C2/N40 ;
    wire \CRT/ssvga_fifo/C2/N35 ;
    wire \CRT/ssvga_fifo/rd_ptr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C103/N20 ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N18 ;
    wire \CRT/ssvga_wbm_if/C1475/N24 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_bc_out[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C26/N18 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C26/N24 ;
    wire \bridge/wishbone_slave_unit/pcim_if_bc_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_bc_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[5]/SRNOT ;
    wire \CRT/ssvga_fifo/C2/N30 ;
    wire \CRT/ssvga_fifo/C2/N25 ;
    wire \CRT/ssvga_fifo/rd_ptr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N30 ;
    wire \CRT/ssvga_wbm_if/C1475/N36 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[7]/SRNOT ;
    wire \CRT/ssvga_fifo/C2/N20 ;
    wire \CRT/ssvga_fifo/C2/N15 ;
    wire \CRT/ssvga_fifo/rd_ptr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N42 ;
    wire \CRT/ssvga_wbm_if/C1475/N48 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[9]/SRNOT ;
    wire \CRT/ssvga_fifo/C2/N10 ;
    wire \CRT/ssvga_fifo/C2/N5 ;
    wire \CRT/ssvga_fifo/rd_ptr[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/FROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/reg_empty ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FFY/SET ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[1]/SRNOT ;
    wire \CRT/ssvga_fifo/C751/N6 ;
    wire \CRT/ssvga_fifo/C751/N11 ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[3]/SRNOT ;
    wire \CRT/ssvga_fifo/C751/N16 ;
    wire \CRT/ssvga_fifo/C751/N21 ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N306 ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N307 ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[3]/FFY/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[3]/FFX/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[5]/SRNOT ;
    wire \CRT/ssvga_fifo/C751/N26 ;
    wire \CRT/ssvga_fifo/C751/N31 ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N308 ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[4]/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[4]/FFY/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[7]/SRNOT ;
    wire \CRT/ssvga_fifo/C751/N36 ;
    wire \CRT/ssvga_fifo/C751/N41 ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N288 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N289 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/SRNOT ;
    wire N12588;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[9]/SRNOT ;
    wire \CRT/ssvga_fifo/C751/N46 ;
    wire \CRT/ssvga_fifo/C751/N51 ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N290 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[0]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[0]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty121 ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[1]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[1]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[2]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[2]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[2]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[0]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C83/N38 ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[0]/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[3]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[3]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_be_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[1]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C83/N27 ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[1]/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[2]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C83/N15 ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[2]/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/c_state[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/inGreyCount[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/inGreyCount[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/inGreyCount[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/inGreyCount[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/inGreyCount[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/delete_status_bit13/SRNOT ;
    wire \bridge/configuration/C384/N3 ;
    wire \bridge/configuration/C383/N3 ;
    wire \bridge/configuration/delete_status_bit13/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/delete_status_bit13/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/SRNOT ;
    wire N12589;
    wire \bridge/wishbone_slave_unit/wishbone_slave/wdel_completion_allow ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/output_backup/mas_ad_en_out/SRNOT ;
    wire \bridge/output_backup/mas_ad_en_out/GROM ;
    wire \bridge/output_backup/mas_ad_en_out/FROM ;
    wire \bridge/output_backup/mas_ad_en_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty116 ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[1]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N6 ;
    wire \CRT/ssvga_wbm_if/C1474/N11 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos_wbw_full_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/reg_full ;
    wire \bridge/wishbone_slave_unit/fifos_wbw_full_out/FROM ;
    wire \bridge/wishbone_slave_unit/fifos_wbw_full_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_write_performed/BYNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_write_performed/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_write_performed/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_write_performed/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[3]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N16 ;
    wire \CRT/ssvga_wbm_if/C1474/N21 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/parchk_sig_serr_out/SRNOT ;
    wire \bridge/parchk_sig_serr_out/GROM ;
    wire \bridge/parchk_sig_serr_out/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[5]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N26 ;
    wire \CRT/ssvga_wbm_if/C1474/N31 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/state_backoff_reg/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/state_backoff_reg/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/N63 ;
    wire \bridge/pci_target_unit/pci_target_sm/state_backoff_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/state_backoff_reg/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_cbe_en_out/SRNOT ;
    wire \bridge/out_bckp_cbe_en_out/GROM ;
    wire \bridge/out_bckp_cbe_en_out/FROM ;
    wire \bridge/out_bckp_cbe_en_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/delete_status_bit15/SRNOT ;
    wire \bridge/configuration/C382/N3 ;
    wire \bridge/configuration/C381/N3 ;
    wire \bridge/configuration/delete_status_bit15/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/delete_status_bit15/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[7]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N36 ;
    wire \CRT/ssvga_wbm_if/C1474/N41 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[9]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N46 ;
    wire \CRT/ssvga_wbm_if/C1474/N51 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/do_master_abort ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/c_state[0]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/C4/N19 ;
    wire \bridge/pci_target_unit/pci_target_sm/c_state[0]/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/c_state[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/c_state[1]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/C4/N11 ;
    wire \bridge/pci_target_unit/pci_target_sm/c_state[1]/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/c_state[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/reg_empty ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[11]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N56 ;
    wire \CRT/ssvga_wbm_if/C1474/N62 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[2]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N6 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[2]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N12 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[3]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[13]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N66 ;
    wire \CRT/ssvga_wbm_if/C1474/N72 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[4]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N18 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[4]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[5]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N24 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[5]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[15]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N76 ;
    wire \CRT/ssvga_wbm_if/C1474/N81 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_pci_drcomp_pending_out/SRNOT ;
    wire N12603;
    wire \bridge/pciu_pci_drcomp_pending_out/FROM ;
    wire \bridge/pciu_pci_drcomp_pending_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[6]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N30 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[6]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[6]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[7]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N36 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[7]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[16]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1474/N87 ;
    wire \CRT/ssvga_wbm_if/vmaddr_r[16]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[8]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N42 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[8]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[8]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[9]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N48 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[9]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_bc_out[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_bc_out[3]/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync_bc_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/req_comp_pending/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C9/N5 ;
    wire \bridge/pci_target_unit/del_sync/req_comp_pending/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C9/N5 ;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_comp_flush_out/SRNOT ;
    wire \bridge/pci_target_unit/fifos/C2/N5 ;
    wire \bridge/pci_target_unit/del_sync_comp_flush_out/FROM ;
    wire \bridge/pci_target_unit/del_sync_comp_flush_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_comp_flush_out/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C93/N5 ;
    wire \bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/N1860 ;
    wire \bridge/wishbone_slave_unit/fifos/N1861 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_almost_full_in ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_ssvga_en/SRNOT ;
    wire \CRT/ssvga_crtc/C531/N5 ;
    wire \CRT/ssvga_fifo/sync_ssvga_en/FROM ;
    wire \CRT/ssvga_fifo/sync_ssvga_en/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_ssvga_en/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/map/SRNOT ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/n_859 ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/map/FROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/map/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[1]/SRNOT ;
    wire \CRT/ssvga_crtc/C531/N10 ;
    wire \CRT/ssvga_crtc/hcntr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[3]/SRNOT ;
    wire \CRT/ssvga_crtc/C531/N15 ;
    wire \CRT/ssvga_crtc/C531/N20 ;
    wire \CRT/ssvga_crtc/hcntr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[5]/SRNOT ;
    wire \CRT/ssvga_crtc/C531/N25 ;
    wire \CRT/ssvga_crtc/C531/N30 ;
    wire \CRT/ssvga_crtc/hcntr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[7]/SRNOT ;
    wire \CRT/ssvga_crtc/C531/N35 ;
    wire \CRT/ssvga_crtc/C531/N40 ;
    wire \CRT/ssvga_crtc/hcntr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[9]/SRNOT ;
    wire \CRT/ssvga_crtc/C531/N45 ;
    wire \CRT/ssvga_crtc/C531/N50 ;
    wire \CRT/ssvga_crtc/hcntr[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/hcntr[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_trdy_en_out/SRNOT ;
    wire \bridge/out_bckp_trdy_en_out/GROM ;
    wire \bridge/out_bckp_trdy_en_out/FROM ;
    wire \bridge/out_bckp_trdy_en_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N54 ;
    wire \CRT/ssvga_wbm_if/C1475/N60 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N114 ;
    wire \CRT/ssvga_wbm_if/C1475/N120 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N66 ;
    wire \CRT/ssvga_wbm_if/C1475/N72 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/SRNOT ;
    wire \bridge/parity_checker/par_cbe_include ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N174 ;
    wire \CRT/ssvga_wbm_if/C1475/N180 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N126 ;
    wire \CRT/ssvga_wbm_if/C1475/N132 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N78 ;
    wire \CRT/ssvga_wbm_if/C1475/N84 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N138 ;
    wire \CRT/ssvga_wbm_if/C1475/N144 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N90 ;
    wire \CRT/ssvga_wbm_if/C1475/N96 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N150 ;
    wire \CRT/ssvga_wbm_if/C1475/N156 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N102 ;
    wire \CRT/ssvga_wbm_if/C1475/N108 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/SRNOT ;
    wire \CRT/ssvga_wbm_if/C1475/N162 ;
    wire \CRT/ssvga_wbm_if/C1475/N168 ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/data_source/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/data_source/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/data_source/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/data_source/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/req_comp_pending_sample/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C8/N6 ;
    wire \bridge/pci_target_unit/del_sync/req_comp_pending_sample/FROM ;
    wire \bridge/pci_target_unit/del_sync/req_comp_pending_sample/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/req_comp_pending_sample/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/parity_checker/perr_sampled/SRNOT ;
    wire \bridge/parity_checker/perr_sampled_in ;
    wire \bridge/parity_checker/perr_sampled/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/delete_status_bit11/SRNOT ;
    wire \bridge/configuration/C386/N3 ;
    wire \bridge/configuration/C385/N3 ;
    wire \bridge/configuration/delete_status_bit11/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/delete_status_bit11/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_empty ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/N1828 ;
    wire \bridge/wishbone_slave_unit/fifos/N1829 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos_pciw_two_left_out/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_two_left_in ;
    wire \bridge/pci_target_unit/fifos_pciw_two_left_out/FROM ;
    wire \bridge/pci_target_unit/fifos_pciw_two_left_out/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/crtc_vblank/SRNOT ;
    wire N12150;
    wire \CRT/crtc_vblank/FROM ;
    wire \CRT/crtc_vblank/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty101 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_almost_empty ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/inGreyCount[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_frame_out/SRNOT ;
    wire \bridge/out_bckp_frame_out/GROM ;
    wire \bridge/out_bckp_frame_out/FROM ;
    wire \bridge/out_bckp_frame_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_empty ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/outGreyCount[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/outGreyCount[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/outGreyCount[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/outGreyCount[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/outGreyCount[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[1]/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[3]/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[4]/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[4]/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_raddr_0[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/drive_blank_reg/SRNOT ;
    wire \CRT/drive_blank_reg160 ;
    wire \CRT/drive_blank_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/last_int ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[0]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N5 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[0]/FROM ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N5 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit10_8[9]/SRNOT ;
    wire \bridge/configuration/wb_err_cs_bit10_8[9]/GROM ;
    wire \bridge/configuration/wb_err_cs_bit10_8[9]/FROM ;
    wire \bridge/configuration/wb_err_cs_bit10_8[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[3]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N15 ;
    wire \bridge/pci_target_unit/del_sync/C1265/N20 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N15 ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N20 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C78/N44 ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/FROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[5]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N25 ;
    wire \bridge/pci_target_unit/del_sync/C1265/N30 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N25 ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N30 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C78/N31 ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/FROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/SRNOT ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C78/N18 ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/FROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[7]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N35 ;
    wire \bridge/pci_target_unit/del_sync/C1265/N40 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N35 ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N40 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[9]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C1265/N45 ;
    wire \bridge/pci_target_unit/del_sync/C1265/N50 ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N45 ;
    wire \bridge/wishbone_slave_unit/del_sync/C25/N50 ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[10]/SRNOT ;
    wire \bridge/out_bckp_ad_out[10]/GROM ;
    wire \bridge/out_bckp_ad_out[10]/FROM ;
    wire \bridge/out_bckp_ad_out[10]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[11]/SRNOT ;
    wire \bridge/out_bckp_ad_out[11]/GROM ;
    wire \bridge/out_bckp_ad_out[11]/FROM ;
    wire \bridge/out_bckp_ad_out[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[20]/SRNOT ;
    wire \bridge/out_bckp_ad_out[20]/GROM ;
    wire \bridge/out_bckp_ad_out[20]/FROM ;
    wire \bridge/out_bckp_ad_out[20]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[12]/SRNOT ;
    wire \bridge/out_bckp_ad_out[12]/GROM ;
    wire \bridge/out_bckp_ad_out[12]/FROM ;
    wire \bridge/out_bckp_ad_out[12]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[21]/SRNOT ;
    wire \bridge/out_bckp_ad_out[21]/GROM ;
    wire \bridge/out_bckp_ad_out[21]/FROM ;
    wire \bridge/out_bckp_ad_out[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[13]/SRNOT ;
    wire \bridge/out_bckp_ad_out[13]/GROM ;
    wire \bridge/out_bckp_ad_out[13]/FROM ;
    wire \bridge/out_bckp_ad_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[30]/SRNOT ;
    wire \bridge/out_bckp_ad_out[30]/GROM ;
    wire \bridge/out_bckp_ad_out[30]/FROM ;
    wire \bridge/out_bckp_ad_out[30]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[22]/SRNOT ;
    wire \bridge/out_bckp_ad_out[22]/GROM ;
    wire \bridge/out_bckp_ad_out[22]/FROM ;
    wire \bridge/out_bckp_ad_out[22]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[14]/SRNOT ;
    wire \bridge/out_bckp_ad_out[14]/GROM ;
    wire \bridge/out_bckp_ad_out[14]/FROM ;
    wire \bridge/out_bckp_ad_out[14]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[31]/SRNOT ;
    wire \bridge/out_bckp_ad_out[31]/GROM ;
    wire \bridge/out_bckp_ad_out[31]/FROM ;
    wire \bridge/out_bckp_ad_out[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[23]/SRNOT ;
    wire \bridge/out_bckp_ad_out[23]/GROM ;
    wire \bridge/out_bckp_ad_out[23]/FROM ;
    wire \bridge/out_bckp_ad_out[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[15]/SRNOT ;
    wire \bridge/out_bckp_ad_out[15]/GROM ;
    wire \bridge/out_bckp_ad_out[15]/FROM ;
    wire \bridge/out_bckp_ad_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[24]/SRNOT ;
    wire \bridge/out_bckp_ad_out[24]/GROM ;
    wire \bridge/out_bckp_ad_out[24]/FROM ;
    wire \bridge/out_bckp_ad_out[24]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[16]/SRNOT ;
    wire \bridge/out_bckp_ad_out[16]/GROM ;
    wire \bridge/out_bckp_ad_out[16]/FROM ;
    wire \bridge/out_bckp_ad_out[16]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[25]/SRNOT ;
    wire \bridge/out_bckp_ad_out[25]/GROM ;
    wire \bridge/out_bckp_ad_out[25]/FROM ;
    wire \bridge/out_bckp_ad_out[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[17]/SRNOT ;
    wire \bridge/out_bckp_ad_out[17]/GROM ;
    wire \bridge/out_bckp_ad_out[17]/FROM ;
    wire \bridge/out_bckp_ad_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[26]/SRNOT ;
    wire \bridge/out_bckp_ad_out[26]/GROM ;
    wire \bridge/out_bckp_ad_out[26]/FROM ;
    wire \bridge/out_bckp_ad_out[26]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[18]/SRNOT ;
    wire \bridge/out_bckp_ad_out[18]/GROM ;
    wire \bridge/out_bckp_ad_out[18]/FROM ;
    wire \bridge/out_bckp_ad_out[18]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_trdy_out/SRNOT ;
    wire \bridge/out_bckp_trdy_out/GROM ;
    wire \bridge/out_bckp_trdy_out/FROM ;
    wire \bridge/out_bckp_trdy_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N318 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N319 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[27]/SRNOT ;
    wire \bridge/out_bckp_ad_out[27]/GROM ;
    wire \bridge/out_bckp_ad_out[27]/FROM ;
    wire \bridge/out_bckp_ad_out[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[19]/SRNOT ;
    wire \bridge/out_bckp_ad_out[19]/GROM ;
    wire \bridge/out_bckp_ad_out[19]/FROM ;
    wire \bridge/out_bckp_ad_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_tar_ad_en_out/SRNOT ;
    wire \bridge/out_bckp_tar_ad_en_out/GROM ;
    wire \bridge/out_bckp_tar_ad_en_out/FROM ;
    wire \bridge/out_bckp_tar_ad_en_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[28]/SRNOT ;
    wire \bridge/out_bckp_ad_out[28]/GROM ;
    wire \bridge/out_bckp_ad_out[28]/FROM ;
    wire \bridge/out_bckp_ad_out[28]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N320 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_ad_out[29]/SRNOT ;
    wire \bridge/out_bckp_ad_out[29]/GROM ;
    wire \bridge/out_bckp_ad_out[29]/FROM ;
    wire \bridge/out_bckp_ad_out[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N321 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[5]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/SRNOT ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/wdel_addr_hit ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/FROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C25/N6 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C25/N12 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C20/N6 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_perr_out/SRNOT ;
    wire \bridge/out_bckp_perr_out/GROM ;
    wire \bridge/out_bckp_perr_out/FROM ;
    wire \bridge/out_bckp_perr_out/FFY/ASYNC_FF_GSR_OR ;
    wire \ACK_I/SRNOT ;
    wire \ACK_I/GROM ;
    wire \ACK_I/FROM ;
    wire \ACK_I/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_comp_req_pending_out/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/C4/N5 ;
    wire \bridge/pci_target_unit/del_sync_comp_req_pending_out/FROM ;
    wire \bridge/pci_target_unit/del_sync_comp_req_pending_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/C4/N5 ;
    wire \bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_read_processing_out/SRNOT ;
    wire N12601;
    wire \bridge/pci_target_unit/pcit_if_read_processing_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_req_req_pending_out/SRNOT ;
    wire N12591;
    wire \bridge/wishbone_slave_unit/del_sync_req_req_pending_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/C2/N5 ;
    wire \bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_progress/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/read_progress ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_progress/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_progress/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[1]/SRNOT ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[3]/SRNOT ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[5]/SRNOT ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[7]/SRNOT ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_clr/SRNOT ;
    wire \bridge/parity_checker/frame_dec2201 ;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_clr/FROM ;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_clr/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[9]/SRNOT ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FROM ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[1]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFX/SET ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/reset_rty_cnt/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/reset_rty_cnt379 ;
    wire \bridge/pci_target_unit/wishbone_master/reset_rty_cnt/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/reset_rty_cnt/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[10]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N54 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[10]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[10]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[11]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N60 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[11]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[20]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N114 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[20]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[20]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[12]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N66 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[12]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[12]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/parity_checker/pci_perr_en_reg/SRNOT ;
    wire \bridge/parity_checker/pci_perr_en_reg/GROM ;
    wire \bridge/parity_checker/perr_en_crit_gen/perr ;
    wire \bridge/parity_checker/pci_perr_en_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/parity_checker/pci_perr_en_reg/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[21]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N120 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[21]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[13]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N72 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[13]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[30]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N174 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[30]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[30]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[22]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N126 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[22]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[22]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[14]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N78 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[14]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[14]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[31]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N180 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[31]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[23]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N132 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[23]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[15]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N84 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[15]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[24]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N138 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[24]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[24]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[16]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N90 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[16]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[16]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[25]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N144 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[25]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[17]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N96 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[17]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[26]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N150 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[26]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[26]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[18]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N102 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[18]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[18]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[27]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N156 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[27]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[19]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N108 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[19]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N6 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[28]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N162 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[28]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[28]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[29]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3276/N168 ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[29]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N18 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N24 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N30 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N36 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/N2000 ;
    wire \bridge/pci_target_unit/fifos/N2001 ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C0/N6 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N42 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N48 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C17/N5 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_bound/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N53 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3277/N12 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/SRNOT ;
    wire \CRT/ssvga_wbm_if/frame_read_in ;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_from_fifo/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/write_to_fifo ;
    wire \bridge/pci_target_unit/pci_target_sm/read_from_fifo ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_from_fifo/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/rd_from_fifo/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[0]/SRNOT ;
    wire \CRT/ssvga_crtc/C532/N5 ;
    wire \CRT/ssvga_crtc/vcntr[0]/FROM ;
    wire \CRT/ssvga_crtc/vcntr[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[1]/SRNOT ;
    wire \CRT/ssvga_crtc/C532/N10 ;
    wire \CRT/ssvga_crtc/vcntr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[3]/SRNOT ;
    wire \CRT/ssvga_crtc/C532/N15 ;
    wire \CRT/ssvga_crtc/C532/N20 ;
    wire \CRT/ssvga_crtc/vcntr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[5]/SRNOT ;
    wire \CRT/ssvga_crtc/C532/N25 ;
    wire \CRT/ssvga_crtc/C532/N30 ;
    wire \CRT/ssvga_crtc/vcntr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[7]/SRNOT ;
    wire \CRT/ssvga_crtc/C532/N35 ;
    wire \CRT/ssvga_crtc/C532/N40 ;
    wire \CRT/ssvga_crtc/vcntr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/write_req_int327 ;
    wire syn22180;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[9]/SRNOT ;
    wire \CRT/ssvga_crtc/C532/N45 ;
    wire \CRT/ssvga_crtc/C532/N50 ;
    wire \CRT/ssvga_crtc/vcntr[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/vcntr[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/go/SRNOT ;
    wire \CRT/C0/N5 ;
    wire \CRT/go/FROM ;
    wire \CRT/go/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[0]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[0]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[1]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[3]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[3]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[5]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[5]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[5]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[1]/SRNOT ;
    wire \CRT/ssvga_fifo/C750/N6 ;
    wire \CRT/ssvga_fifo/C750/N11 ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/out_bckp_devsel_out/SRNOT ;
    wire \bridge/out_bckp_devsel_out/GROM ;
    wire \bridge/out_bckp_devsel_out/FROM ;
    wire \bridge/out_bckp_devsel_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[7]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[7]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[7]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr[1]/SRNOT ;
    wire \CRT/ssvga_fifo/C0/N40 ;
    wire \CRT/ssvga_fifo/C0/N35 ;
    wire \CRT/ssvga_fifo/wr_ptr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[11]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[11]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[11]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[3]/SRNOT ;
    wire \CRT/ssvga_fifo/C750/N16 ;
    wire \CRT/ssvga_fifo/C750/N21 ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[9]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[9]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[9]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr[3]/SRNOT ;
    wire \CRT/ssvga_fifo/C0/N30 ;
    wire \CRT/ssvga_fifo/C0/N25 ;
    wire \CRT/ssvga_fifo/wr_ptr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[21]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[21]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[21]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[13]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[13]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[13]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[5]/SRNOT ;
    wire \CRT/ssvga_fifo/C750/N26 ;
    wire \CRT/ssvga_fifo/C750/N31 ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N132 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N126 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr[5]/SRNOT ;
    wire \CRT/ssvga_fifo/C0/N20 ;
    wire \CRT/ssvga_fifo/C0/N15 ;
    wire \CRT/ssvga_fifo/wr_ptr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[31]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[31]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[31]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[23]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[23]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[23]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[15]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[15]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[15]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[7]/SRNOT ;
    wire \CRT/ssvga_fifo/C750/N36 ;
    wire \CRT/ssvga_fifo/C750/N41 ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N72 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N66 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N120 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N114 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr[7]/SRNOT ;
    wire \CRT/ssvga_fifo/C0/N10 ;
    wire \CRT/ssvga_fifo/C0/N5 ;
    wire \CRT/ssvga_fifo/wr_ptr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/wr_ptr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w/FROM ;
    wire \syn17012/GROM ;
    wire \syn17012/FROM ;
    wire \syn19385/GROM ;
    wire \syn19385/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/stop_w/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/stop_w/FROM ;
    wire \syn17093/GROM ;
    wire \syn17093/FROM ;
    wire \syn179249/GROM ;
    wire \syn179249/FROM ;
    wire \SDAT_O[31]/GROM ;
    wire \SDAT_O[31]/FROM ;
    wire \syn177518/GROM ;
    wire \syn177518/FROM ;
    wire \syn177514/GROM ;
    wire \syn177514/FROM ;
    wire \bridge/configuration/C2308/GROM ;
    wire \bridge/configuration/C2308/FROM ;
    wire \syn177396/GROM ;
    wire \syn177396/FROM ;
    wire \syn177397/GROM ;
    wire \syn177397/FROM ;
    wire \syn17813/GROM ;
    wire \syn17813/FROM ;
    wire \bridge/configuration/C2370/GROM ;
    wire \bridge/configuration/C2370/FROM ;
    wire \bridge/configuration/C2338/GROM ;
    wire \bridge/configuration/C2338/FROM ;
    wire \bridge/configuration/C2354/GROM ;
    wire \bridge/configuration/C2354/FROM ;
    wire \bridge/configuration/C2340/GROM ;
    wire \bridge/configuration/C2340/FROM ;
    wire \syn177519/GROM ;
    wire \syn177519/FROM ;
    wire \bridge/configuration/C2356/GROM ;
    wire \bridge/configuration/C2356/FROM ;
    wire \syn120377/GROM ;
    wire \syn120377/FROM ;
    wire \syn177508/GROM ;
    wire \syn177508/FROM ;
    wire \bridge/configuration/C2322/GROM ;
    wire \bridge/configuration/C2322/FROM ;
    wire \syn177509/GROM ;
    wire \syn177509/FROM ;
    wire \bridge/configuration/C2302/GROM ;
    wire \bridge/configuration/C2302/FROM ;
    wire \syn177512/GROM ;
    wire \syn177512/FROM ;
    wire \bridge/configuration/C2368/GROM ;
    wire \bridge/configuration/C2368/FROM ;
    wire \bridge/configuration/C2360/GROM ;
    wire \bridge/configuration/C2360/FROM ;
    wire \bridge/configuration/C2320/GROM ;
    wire \bridge/configuration/C2320/FROM ;
    wire \syn17836/GROM ;
    wire \syn17836/FROM ;
    wire \syn177416/GROM ;
    wire \syn177416/FROM ;
    wire \syn24326/GROM ;
    wire \syn24326/FROM ;
    wire \syn24559/GROM ;
    wire \syn24559/FROM ;
    wire \syn177532/GROM ;
    wire \syn177532/FROM ;
    wire \SDAT_O[30]/GROM ;
    wire \SDAT_O[30]/FROM ;
    wire \syn177580/GROM ;
    wire \syn177580/FROM ;
    wire \bridge/configuration/C2304/GROM ;
    wire \bridge/configuration/C2304/FROM ;
    wire \syn177581/GROM ;
    wire \syn177581/FROM ;
    wire \syn177573/GROM ;
    wire \syn177573/FROM ;
    wire \syn16917/GROM ;
    wire \syn16917/FROM ;
    wire \SDAT_O[29]/GROM ;
    wire \SDAT_O[29]/FROM ;
    wire \syn177616/GROM ;
    wire \syn177616/FROM ;
    wire \bridge/configuration/C2318/GROM ;
    wire \bridge/configuration/C2318/FROM ;
    wire \syn177620/GROM ;
    wire \syn177620/FROM ;
    wire \SDAT_O[28]/GROM ;
    wire \SDAT_O[28]/FROM ;
    wire \syn177664/GROM ;
    wire \syn177664/FROM ;
    wire \syn177665/GROM ;
    wire \syn177665/FROM ;
    wire \syn177669/GROM ;
    wire \syn177669/FROM ;
    wire \SDAT_O[27]/GROM ;
    wire \SDAT_O[27]/FROM ;
    wire \syn50278/GROM ;
    wire \syn50278/FROM ;
    wire \syn177703/GROM ;
    wire \syn177703/FROM ;
    wire \syn177704/GROM ;
    wire \syn177704/FROM ;
    wire \syn177701/GROM ;
    wire \syn177701/FROM ;
    wire \SDAT_O[26]/GROM ;
    wire \SDAT_O[26]/FROM ;
    wire \syn177743/GROM ;
    wire \syn177743/FROM ;
    wire \syn177734/GROM ;
    wire \syn177734/FROM ;
    wire \syn177744/GROM ;
    wire \syn177744/FROM ;
    wire \SDAT_O[25]/GROM ;
    wire \SDAT_O[25]/FROM ;
    wire \syn50276/GROM ;
    wire \syn50276/FROM ;
    wire \syn177782/GROM ;
    wire \syn177782/FROM ;
    wire \SDAT_O[24]/GROM ;
    wire \SDAT_O[24]/FROM ;
    wire \syn177822/GROM ;
    wire \syn177822/FROM ;
    wire \syn177826/GROM ;
    wire \syn177826/FROM ;
    wire \SDAT_O[23]/GROM ;
    wire \SDAT_O[23]/FROM ;
    wire \syn177864/GROM ;
    wire \syn177864/FROM ;
    wire \syn177865/GROM ;
    wire \syn177865/FROM ;
    wire \syn177855/GROM ;
    wire \syn177855/FROM ;
    wire \syn177858/GROM ;
    wire \syn177858/FROM ;
    wire \bridge/configuration/C2296/GROM ;
    wire \bridge/configuration/C2296/FROM ;
    wire \SDAT_O[22]/GROM ;
    wire \SDAT_O[22]/FROM ;
    wire \syn177897/GROM ;
    wire \syn177897/FROM ;
    wire \syn177898/GROM ;
    wire \syn177898/FROM ;
    wire \syn177888/GROM ;
    wire \syn177888/FROM ;
    wire \syn177891/GROM ;
    wire \syn177891/FROM ;
    wire \SDAT_O[21]/GROM ;
    wire \SDAT_O[21]/FROM ;
    wire \syn177927/GROM ;
    wire \syn177927/FROM ;
    wire \syn177931/GROM ;
    wire \syn177931/FROM ;
    wire \syn177936/GROM ;
    wire \syn177936/FROM ;
    wire \SDAT_O[20]/GROM ;
    wire \SDAT_O[20]/FROM ;
    wire \syn177960/GROM ;
    wire \syn177960/FROM ;
    wire \syn177964/GROM ;
    wire \syn177964/FROM ;
    wire \syn177969/GROM ;
    wire \syn177969/FROM ;
    wire \SDAT_O[19]/GROM ;
    wire \SDAT_O[19]/FROM ;
    wire \syn177997/GROM ;
    wire \syn177997/FROM ;
    wire \syn177998/GROM ;
    wire \syn177998/FROM ;
    wire \syn177988/GROM ;
    wire \syn177988/FROM ;
    wire \syn177991/GROM ;
    wire \syn177991/FROM ;
    wire \SDAT_O[18]/GROM ;
    wire \SDAT_O[18]/FROM ;
    wire \syn178030/GROM ;
    wire \syn178030/FROM ;
    wire \syn178031/GROM ;
    wire \syn178031/FROM ;
    wire \syn178021/GROM ;
    wire \syn178021/FROM ;
    wire \syn178024/GROM ;
    wire \syn178024/FROM ;
    wire \SDAT_O[17]/GROM ;
    wire \SDAT_O[17]/FROM ;
    wire \syn178060/GROM ;
    wire \syn178060/FROM ;
    wire \syn178064/GROM ;
    wire \syn178064/FROM ;
    wire \syn178069/GROM ;
    wire \syn178069/FROM ;
    wire \SDAT_O[16]/GROM ;
    wire \SDAT_O[16]/FROM ;
    wire \syn178101/GROM ;
    wire \syn178101/FROM ;
    wire \syn178102/GROM ;
    wire \syn178102/FROM ;
    wire \syn17772/GROM ;
    wire \syn17772/FROM ;
    wire \SDAT_O[15]/GROM ;
    wire \SDAT_O[15]/FROM ;
    wire \syn178139/GROM ;
    wire \syn178139/FROM ;
    wire \syn178140/GROM ;
    wire \syn178140/FROM ;
    wire \syn178130/GROM ;
    wire \syn178130/FROM ;
    wire \syn178133/GROM ;
    wire \syn178133/FROM ;
    wire \syn178144/GROM ;
    wire \syn178144/FROM ;
    wire \SDAT_O[14]/GROM ;
    wire \SDAT_O[14]/FROM ;
    wire \syn178174/GROM ;
    wire \syn178174/FROM ;
    wire \syn178175/GROM ;
    wire \syn178175/FROM ;
    wire \syn178165/GROM ;
    wire \syn178165/FROM ;
    wire \syn178168/GROM ;
    wire \syn178168/FROM ;
    wire \SDAT_O[13]/GROM ;
    wire \SDAT_O[13]/FROM ;
    wire \syn18511/GROM ;
    wire \syn18511/FROM ;
    wire \syn178206/GROM ;
    wire \syn178206/FROM ;
    wire \syn178208/GROM ;
    wire \syn178208/FROM ;
    wire \syn178213/GROM ;
    wire \syn178213/FROM ;
    wire \SDAT_O[12]/GROM ;
    wire \SDAT_O[12]/FROM ;
    wire \syn178245/GROM ;
    wire \syn178245/FROM ;
    wire \syn178246/GROM ;
    wire \syn178246/FROM ;
    wire \SDAT_O[11]/GROM ;
    wire \SDAT_O[11]/FROM ;
    wire \syn178265/GROM ;
    wire \syn178265/FROM ;
    wire \syn178266/GROM ;
    wire \syn178266/FROM ;
    wire \SDAT_O[10]/GROM ;
    wire \SDAT_O[10]/FROM ;
    wire \syn178294/GROM ;
    wire \syn178294/FROM ;
    wire \syn16936/GROM ;
    wire \syn16936/FROM ;
    wire \syn178292/GROM ;
    wire \syn178292/FROM ;
    wire \SDAT_O[9]/GROM ;
    wire \SDAT_O[9]/FROM ;
    wire \syn178312/GROM ;
    wire \syn178312/FROM ;
    wire \SDAT_O[8]/GROM ;
    wire \SDAT_O[8]/FROM ;
    wire \syn178340/GROM ;
    wire \syn178340/FROM ;
    wire \syn178341/GROM ;
    wire \syn178341/FROM ;
    wire \syn178334/GROM ;
    wire \syn178334/FROM ;
    wire \syn178338/GROM ;
    wire \syn178338/FROM ;
    wire \SDAT_O[7]/GROM ;
    wire \SDAT_O[7]/FROM ;
    wire \syn178357/GROM ;
    wire \syn178357/FROM ;
    wire \SDAT_O[6]/GROM ;
    wire \SDAT_O[6]/FROM ;
    wire \syn178375/GROM ;
    wire \syn178375/FROM ;
    wire \SDAT_O[5]/GROM ;
    wire \SDAT_O[5]/FROM ;
    wire \syn178393/GROM ;
    wire \syn178393/FROM ;
    wire \syn178392/GROM ;
    wire \syn178392/FROM ;
    wire \SDAT_O[4]/GROM ;
    wire \SDAT_O[4]/FROM ;
    wire \syn178410/GROM ;
    wire \syn178410/FROM ;
    wire \SDAT_O[3]/GROM ;
    wire \SDAT_O[3]/FROM ;
    wire \syn178435/GROM ;
    wire \syn178435/FROM ;
    wire \syn178432/GROM ;
    wire \syn178432/FROM ;
    wire \SDAT_O[2]/GROM ;
    wire \SDAT_O[2]/FROM ;
    wire \syn18765/GROM ;
    wire \syn18765/FROM ;
    wire \syn178459/GROM ;
    wire \syn178459/FROM ;
    wire \syn178449/GROM ;
    wire \syn178449/FROM ;
    wire \SDAT_O[1]/GROM ;
    wire \SDAT_O[1]/FROM ;
    wire \syn178488/GROM ;
    wire \syn178488/FROM ;
    wire \syn178489/GROM ;
    wire \syn178489/FROM ;
    wire \SDAT_O[0]/GROM ;
    wire \SDAT_O[0]/FROM ;
    wire \syn178523/GROM ;
    wire \syn178523/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N35/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N35/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow/FROM ;
    wire \syn16935/GROM ;
    wire \syn16935/FROM ;
    wire \CRT/ssvga_wbm_if/S_41/cell0/GROM ;
    wire \CRT/ssvga_wbm_if/S_41/cell0/FROM ;
    wire \syn177319/GROM ;
    wire \syn177319/FROM ;
    wire \syn177320/GROM ;
    wire \syn177320/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N30/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N30/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N24/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N24/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N18/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N18/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N12/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N12/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N6/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C6/N6/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_rallow/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_rallow/FROM ;
    wire \bridge/pci_target_unit/fifos/C9/N30/GROM ;
    wire \bridge/pci_target_unit/fifos/C9/N30/FROM ;
    wire \bridge/pci_target_unit/fifos/C9/N24/GROM ;
    wire \bridge/pci_target_unit/fifos/C9/N24/FROM ;
    wire \bridge/pci_target_unit/fifos/C9/N18/GROM ;
    wire \bridge/pci_target_unit/fifos/C9/N18/FROM ;
    wire \bridge/pci_target_unit/fifos/C9/N12/GROM ;
    wire \bridge/pci_target_unit/fifos/C9/N12/FROM ;
    wire \bridge/pci_target_unit/fifos/C9/N6/GROM ;
    wire \bridge/pci_target_unit/fifos/C9/N6/FROM ;
    wire \syn179246/GROM ;
    wire \syn179246/FROM ;
    wire \syn179247/GROM ;
    wire \syn179247/FROM ;
    wire \syn179248/GROM ;
    wire \syn179248/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy/FROM ;
    wire \syn179287/GROM ;
    wire \syn179287/FROM ;
    wire \syn19968/GROM ;
    wire \syn19968/FROM ;
    wire \CRT/fifo_wr_en/GROM ;
    wire \CRT/fifo_wr_en/FROM ;
    wire \syn17116/GROM ;
    wire \syn17116/FROM ;
    wire \syn16914/GROM ;
    wire \syn16914/FROM ;
    wire \syn179881/GROM ;
    wire \syn179881/FROM ;
    wire \syn20662/GROM ;
    wire \syn20662/FROM ;
    wire \syn180051/GROM ;
    wire \syn180051/FROM ;
    wire \bridge/configuration/C1929/GROM ;
    wire \bridge/configuration/C1929/FROM ;
    wire \syn180183/GROM ;
    wire \syn180183/FROM ;
    wire \syn20739/GROM ;
    wire \syn20739/FROM ;
    wire \syn17015/GROM ;
    wire \syn17015/FROM ;
    wire \syn17014/GROM ;
    wire \syn17014/FROM ;
    wire \syn16985/GROM ;
    wire \syn16985/FROM ;
    wire \syn180247/GROM ;
    wire \syn180247/FROM ;
    wire \syn180240/GROM ;
    wire \syn180240/FROM ;
    wire \syn180248/GROM ;
    wire \syn180248/FROM ;
    wire \syn20947/GROM ;
    wire \syn20947/FROM ;
    wire \syn180417/GROM ;
    wire \syn180417/FROM ;
    wire \bridge/configuration/C1989/GROM ;
    wire \bridge/configuration/C1989/FROM ;
    wire \syn180418/GROM ;
    wire \syn180418/FROM ;
    wire \bridge/configuration/C1971/GROM ;
    wire \bridge/configuration/C1971/FROM ;
    wire \syn180440/GROM ;
    wire \syn180440/FROM ;
    wire \syn16929/GROM ;
    wire \syn16929/FROM ;
    wire \syn20987/GROM ;
    wire \syn20987/FROM ;
    wire \syn180490/GROM ;
    wire \syn180490/FROM ;
    wire \syn180535/GROM ;
    wire \syn180535/FROM ;
    wire \syn16927/GROM ;
    wire \syn16927/FROM ;
    wire \syn180582/GROM ;
    wire \syn180582/FROM ;
    wire \syn180580/GROM ;
    wire \syn180580/FROM ;
    wire \syn136384/GROM ;
    wire \syn136384/FROM ;
    wire \syn21143/GROM ;
    wire \syn21143/FROM ;
    wire \syn180672/GROM ;
    wire \syn180672/FROM ;
    wire \syn180719/GROM ;
    wire \syn180719/FROM ;
    wire \syn180765/GROM ;
    wire \syn180765/FROM ;
    wire \syn21298/GROM ;
    wire \syn21298/FROM ;
    wire \syn180855/GROM ;
    wire \syn180855/FROM ;
    wire \syn21430/GROM ;
    wire \syn21430/FROM ;
    wire \syn181000/GROM ;
    wire \syn181000/FROM ;
    wire \syn181001/GROM ;
    wire \syn181001/FROM ;
    wire \syn21407/GROM ;
    wire \syn21407/FROM ;
    wire \bridge/configuration/C1953/GROM ;
    wire \bridge/configuration/C1953/FROM ;
    wire \syn181008/GROM ;
    wire \syn181008/FROM ;
    wire \syn21585/GROM ;
    wire \syn21585/FROM ;
    wire \syn181201/GROM ;
    wire \syn181201/FROM ;
    wire \syn181217/GROM ;
    wire \syn181217/FROM ;
    wire \syn21625/GROM ;
    wire \syn21625/FROM ;
    wire \syn181272/GROM ;
    wire \syn181272/FROM ;
    wire \syn181520/GROM ;
    wire \syn181520/FROM ;
    wire \syn181498/GROM ;
    wire \syn181498/FROM ;
    wire \syn181499/GROM ;
    wire \syn181499/FROM ;
    wire \syn181497/GROM ;
    wire \syn181497/FROM ;
    wire \syn181521/GROM ;
    wire \syn181521/FROM ;
    wire \syn181500/GROM ;
    wire \syn181500/FROM ;
    wire \syn181501/GROM ;
    wire \syn181501/FROM ;
    wire \syn181502/GROM ;
    wire \syn181502/FROM ;
    wire \syn181522/GROM ;
    wire \syn181522/FROM ;
    wire \syn181504/GROM ;
    wire \syn181504/FROM ;
    wire \syn181505/GROM ;
    wire \syn181505/FROM ;
    wire \syn181506/GROM ;
    wire \syn181506/FROM ;
    wire \syn181508/GROM ;
    wire \syn181508/FROM ;
    wire \syn181510/GROM ;
    wire \syn181510/FROM ;
    wire \N12544/GROM ;
    wire \N12544/FROM ;
    wire \bridge/pci_target_unit/pcit_sm_load_medium_reg_out/GROM ;
    wire \bridge/pci_target_unit/pcit_sm_load_medium_reg_out/FROM ;
    wire \syn18863/GROM ;
    wire \syn18863/FROM ;
    wire \syn18858/GROM ;
    wire \syn18858/FROM ;
    wire \syn17669/GROM ;
    wire \syn17669/FROM ;
    wire \syn177570/GROM ;
    wire \syn177570/FROM ;
    wire \syn177658/GROM ;
    wire \syn177658/FROM ;
    wire \syn177781/GROM ;
    wire \syn177781/FROM ;
    wire \syn177924/GROM ;
    wire \syn177924/FROM ;
    wire \syn177957/GROM ;
    wire \syn177957/FROM ;
    wire \syn178057/GROM ;
    wire \syn178057/FROM ;
    wire \syn178095/GROM ;
    wire \syn178095/FROM ;
    wire \syn178239/GROM ;
    wire \syn178239/FROM ;
    wire \syn178522/GROM ;
    wire \syn178522/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N30/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N30/FROM ;
    wire \syn17087/GROM ;
    wire \syn17087/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/cell8/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/cell8/FROM ;
    wire \syn17086/GROM ;
    wire \syn17086/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N24/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N24/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N18/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N18/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N12/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N12/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N6/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N6/FROM ;
    wire \syn19397/GROM ;
    wire \syn19397/FROM ;
    wire \bridge/pci_target_unit/fifos/C10/N30/GROM ;
    wire \bridge/pci_target_unit/fifos/C10/N30/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[1]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[1]/FROM ;
    wire \bridge/pci_target_unit/fifos/C10/N24/GROM ;
    wire \bridge/pci_target_unit/fifos/C10/N24/FROM ;
    wire \bridge/pci_target_unit/fifos/C10/N18/GROM ;
    wire \bridge/pci_target_unit/fifos/C10/N18/FROM ;
    wire \bridge/pci_target_unit/fifos/C10/N12/GROM ;
    wire \bridge/pci_target_unit/fifos/C10/N12/FROM ;
    wire \bridge/pci_target_unit/fifos/C10/N6/GROM ;
    wire \bridge/pci_target_unit/fifos/C10/N6/FROM ;
    wire \bridge/pci_target_unit/fifos/in_count_en/GROM ;
    wire \bridge/pci_target_unit/fifos/in_count_en/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w_frm/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w_frm/FROM ;
    wire \bridge/configuration/C285/N34/GROM ;
    wire \bridge/configuration/C285/N34/FROM ;
    wire \syn20406/GROM ;
    wire \syn20406/FROM ;
    wire \syn20371/GROM ;
    wire \syn20371/FROM ;
    wire \syn179694/GROM ;
    wire \syn179694/FROM ;
    wire \syn179711/GROM ;
    wire \syn179711/FROM ;
    wire \syn179707/GROM ;
    wire \syn179707/FROM ;
    wire \bridge/configuration/C1959/GROM ;
    wire \bridge/configuration/C1959/FROM ;
    wire \syn179709/GROM ;
    wire \syn179709/FROM ;
    wire \syn20486/GROM ;
    wire \syn20486/FROM ;
    wire \syn179855/GROM ;
    wire \syn179855/FROM ;
    wire \syn179846/GROM ;
    wire \syn179846/FROM ;
    wire \syn20502/GROM ;
    wire \syn20502/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C155/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C155/FROM ;
    wire \syn179882/GROM ;
    wire \syn179882/FROM ;
    wire \bridge/output_backup/data_load/GROM ;
    wire \bridge/output_backup/data_load/FROM ;
    wire \syn20532/GROM ;
    wire \syn20532/FROM ;
    wire \syn20523/GROM ;
    wire \syn20523/FROM ;
    wire \syn179919/GROM ;
    wire \syn179919/FROM ;
    wire \syn20564/GROM ;
    wire \syn20564/FROM ;
    wire \syn179960/GROM ;
    wire \syn179960/FROM ;
    wire \syn20598/GROM ;
    wire \syn20598/FROM ;
    wire \syn20611/GROM ;
    wire \syn20611/FROM ;
    wire \syn20635/GROM ;
    wire \syn20635/FROM ;
    wire \syn180031/GROM ;
    wire \syn180031/FROM ;
    wire \syn17110/GROM ;
    wire \syn17110/FROM ;
    wire \syn180032/GROM ;
    wire \syn180032/FROM ;
    wire \syn20672/GROM ;
    wire \syn20672/FROM ;
    wire \syn20688/GROM ;
    wire \syn20688/FROM ;
    wire \syn180082/GROM ;
    wire \syn180082/FROM ;
    wire \syn20701/GROM ;
    wire \syn20701/FROM ;
    wire \syn20720/GROM ;
    wire \syn20720/FROM ;
    wire \syn20759/GROM ;
    wire \syn20759/FROM ;
    wire \syn180176/GROM ;
    wire \syn180176/FROM ;
    wire \syn137911/GROM ;
    wire \syn137911/FROM ;
    wire \syn180212/GROM ;
    wire \syn180212/FROM ;
    wire \syn20817/GROM ;
    wire \syn20817/FROM ;
    wire \syn20835/GROM ;
    wire \syn20835/FROM ;
    wire \syn180282/GROM ;
    wire \syn180282/FROM ;
    wire \syn180321/GROM ;
    wire \syn180321/FROM ;
    wire \syn180322/GROM ;
    wire \syn180322/FROM ;
    wire \syn20882/GROM ;
    wire \syn20882/FROM ;
    wire \syn180373/GROM ;
    wire \syn180373/FROM ;
    wire \syn180374/GROM ;
    wire \syn180374/FROM ;
    wire \syn20922/GROM ;
    wire \syn20922/FROM ;
    wire \syn180387/GROM ;
    wire \syn180387/FROM ;
    wire \syn20963/GROM ;
    wire \syn20963/FROM ;
    wire \syn21003/GROM ;
    wire \syn21003/FROM ;
    wire \syn180528/GROM ;
    wire \syn180528/FROM ;
    wire \syn180529/GROM ;
    wire \syn180529/FROM ;
    wire \syn21041/GROM ;
    wire \syn21041/FROM ;
    wire \syn21080/GROM ;
    wire \syn21080/FROM ;
    wire \syn180569/GROM ;
    wire \syn180569/FROM ;
    wire \syn180570/GROM ;
    wire \syn180570/FROM ;
    wire \syn21104/GROM ;
    wire \syn21104/FROM ;
    wire \syn180628/GROM ;
    wire \syn180628/FROM ;
    wire \syn21158/GROM ;
    wire \syn21158/FROM ;
    wire \syn21197/GROM ;
    wire \syn21197/FROM ;
    wire \syn180706/GROM ;
    wire \syn180706/FROM ;
    wire \syn180707/GROM ;
    wire \syn180707/FROM ;
    wire \syn21235/GROM ;
    wire \syn21235/FROM ;
    wire \syn180752/GROM ;
    wire \syn180752/FROM ;
    wire \syn180753/GROM ;
    wire \syn180753/FROM ;
    wire \syn21259/GROM ;
    wire \syn21259/FROM ;
    wire \syn180811/GROM ;
    wire \syn180811/FROM ;
    wire \syn21313/GROM ;
    wire \syn21313/FROM ;
    wire \syn21346/GROM ;
    wire \syn21346/FROM ;
    wire \syn180888/GROM ;
    wire \syn180888/FROM ;
    wire \syn180906/GROM ;
    wire \syn180906/FROM ;
    wire \syn21385/GROM ;
    wire \syn21385/FROM ;
    wire \syn180940/GROM ;
    wire \syn180940/FROM ;
    wire \syn180961/GROM ;
    wire \syn180961/FROM ;
    wire \syn21462/GROM ;
    wire \syn21462/FROM ;
    wire \syn181045/GROM ;
    wire \syn181045/FROM ;
    wire \syn21479/GROM ;
    wire \syn21479/FROM ;
    wire \syn181062/GROM ;
    wire \syn181062/FROM ;
    wire \syn21465/GROM ;
    wire \syn21465/FROM ;
    wire \syn120365/GROM ;
    wire \syn120365/FROM ;
    wire \syn21511/GROM ;
    wire \syn21511/FROM ;
    wire \syn181096/GROM ;
    wire \syn181096/FROM ;
    wire \syn181114/GROM ;
    wire \syn181114/FROM ;
    wire \syn21552/GROM ;
    wire \syn21552/FROM ;
    wire \syn181147/GROM ;
    wire \syn181147/FROM ;
    wire \syn181165/GROM ;
    wire \syn181165/FROM ;
    wire \syn21601/GROM ;
    wire \syn21601/FROM ;
    wire \syn21641/GROM ;
    wire \syn21641/FROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C749/GROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C749/FROM ;
    wire \syn181511/GROM ;
    wire \syn181511/FROM ;
    wire \syn22093/GROM ;
    wire \syn22093/FROM ;
    wire \syn22083/GROM ;
    wire \syn22083/FROM ;
    wire \N12382/GROM ;
    wire \N12382/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/C81/N3/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/C81/N3/FROM ;
    wire \syn17011/GROM ;
    wire \syn17011/FROM ;
    wire \N12543/GROM ;
    wire \N12543/FROM ;
    wire \syn22771/GROM ;
    wire \syn22771/FROM ;
    wire \syn19709/GROM ;
    wire \syn19709/FROM ;
    wire \syn179112/GROM ;
    wire \syn179112/FROM ;
    wire \syn179113/GROM ;
    wire \syn179113/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/change_state/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/change_state/FROM ;
    wire \CRT/ssvga_fifo/S_28/cell0/GROM ;
    wire \CRT/ssvga_fifo/S_28/cell0/FROM ;
    wire \syn177262/GROM ;
    wire \syn177262/FROM ;
    wire \syn177263/GROM ;
    wire \syn177263/FROM ;
    wire \syn177264/GROM ;
    wire \syn177264/FROM ;
    wire \CRT/ssvga_fifo/C6/N54/GROM ;
    wire \CRT/ssvga_fifo/C6/N54/FROM ;
    wire \syn17811/GROM ;
    wire \syn17811/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/devs_w_frm/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/devs_w_frm/FROM ;
    wire \syn20373/GROM ;
    wire \syn20373/FROM ;
    wire \syn179986/GROM ;
    wire \syn179986/FROM ;
    wire \syn180030/GROM ;
    wire \syn180030/FROM ;
    wire \syn180120/GROM ;
    wire \syn180120/FROM ;
    wire \syn180180/GROM ;
    wire \syn180180/FROM ;
    wire \syn180198/GROM ;
    wire \syn180198/FROM ;
    wire \syn181113/GROM ;
    wire \syn181113/FROM ;
    wire \N12383/GROM ;
    wire \N12383/FROM ;
    wire \syn181563/GROM ;
    wire \syn181563/FROM ;
    wire \N12033/GROM ;
    wire \N12033/FROM ;
    wire \bridge/parity_checker/non_critical_par/GROM ;
    wire \bridge/parity_checker/non_critical_par/FROM ;
    wire \bridge/parity_checker/syn3156/GROM ;
    wire \bridge/parity_checker/syn3156/FROM ;
    wire \syn177213/GROM ;
    wire \syn177213/FROM ;
    wire \syn18066/GROM ;
    wire \syn18066/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N33/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/C3/N33/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135/FROM ;
    wire \syn178898/GROM ;
    wire \syn178898/FROM ;
    wire \syn19590/GROM ;
    wire \syn19590/FROM ;
    wire \N12510/GROM ;
    wire \N12510/FROM ;
    wire \syn179261/GROM ;
    wire \syn179261/FROM ;
    wire \syn179382/GROM ;
    wire \syn179382/FROM ;
    wire \syn16986/GROM ;
    wire \syn16986/FROM ;
    wire \syn179572/GROM ;
    wire \syn179572/FROM ;
    wire \N12237/GROM ;
    wire \N12237/FROM ;
    wire \bridge/configuration/C281/N3/GROM ;
    wire \bridge/configuration/C281/N3/FROM ;
    wire \syn180181/GROM ;
    wire \syn180181/FROM ;
    wire \syn181624/GROM ;
    wire \syn181624/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/data_be_load/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/data_be_load/FROM ;
    wire \syn182015/GROM ;
    wire \syn182015/FROM ;
    wire \syn182018/GROM ;
    wire \syn182018/FROM ;
    wire \syn22805/GROM ;
    wire \syn22805/FROM ;
    wire \syn17006/GROM ;
    wire \syn17006/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame/FROM ;
    wire \syn177380/GROM ;
    wire \syn177380/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy/FROM ;
    wire \N12151/GROM ;
    wire \N12151/FROM ;
    wire \bridge/configuration/C343/N5/GROM ;
    wire \bridge/configuration/C343/N5/FROM ;
    wire \bridge/configuration/C289/N9/GROM ;
    wire \bridge/configuration/C289/N9/FROM ;
    wire \syn182016/GROM ;
    wire \syn182016/FROM ;
    wire \syn182017/GROM ;
    wire \syn182017/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_clear/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_clear/FROM ;
    wire \syn23022/GROM ;
    wire \syn23022/FROM ;
    wire \syn182406/GROM ;
    wire \syn182406/FROM ;
    wire \syn23263/GROM ;
    wire \syn23263/FROM ;
    wire \syn182488/GROM ;
    wire \syn182488/FROM ;
    wire \syn182538/GROM ;
    wire \syn182538/FROM ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0/FROM ;
    wire \syn23568/GROM ;
    wire \syn23568/FROM ;
    wire \syn182579/GROM ;
    wire \syn182579/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0/FROM ;
    wire \bridge/parity_checker/data_par/GROM ;
    wire \bridge/parity_checker/data_par/FROM ;
    wire \bridge/parity_checker/syn3204/GROM ;
    wire \bridge/parity_checker/syn3204/FROM ;
    wire \bridge/wishbone_slave_unit/wbs_sm_cbe_out[3]/GROM ;
    wire \bridge/wishbone_slave_unit/wbs_sm_cbe_out[3]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_control_out[1]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_control_out[1]/FROM ;
    wire \N12164/GROM ;
    wire \N12164/FROM ;
    wire \bridge/pci_mux_irdy_in/GROM ;
    wire \bridge/pci_mux_irdy_in/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync_burst_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_burst_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[4]/FFY/SET ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/trdy_asserted_reg/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/trdy_asserted_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/req_done_reg/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/req_done_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[12]/SRNOT ;
    wire \bridge/configuration/config_addr[12]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[12]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[22]/SRNOT ;
    wire \bridge/configuration/config_addr[22]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[22]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[14]/SRNOT ;
    wire \bridge/configuration/config_addr[14]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[14]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[23]/SRNOT ;
    wire \bridge/configuration/config_addr[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[15]/SRNOT ;
    wire \bridge/configuration/config_addr[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[16]/SRNOT ;
    wire \bridge/configuration/config_addr[16]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[18]/SRNOT ;
    wire \bridge/configuration/config_addr[18]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[18]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[21]/SRNOT ;
    wire \bridge/configuration/pci_addr_mask1[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[13]/SRNOT ;
    wire \bridge/configuration/pci_addr_mask1[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[20]/SRNOT ;
    wire \bridge/configuration/config_addr[20]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[20]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_bc_out[1]/SRNOT ;
    wire \bridge/pciu_err_bc_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_bc_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_am1_out[19]/SRNOT ;
    wire \bridge/conf_pci_am1_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_am1_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[23]/SRNOT ;
    wire \bridge/configuration/pci_addr_mask1[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[15]/SRNOT ;
    wire \bridge/configuration/pci_addr_mask1[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_bc_out[3]/SRNOT ;
    wire \bridge/pciu_err_bc_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_err_bc_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_am1_out[13]/SRNOT ;
    wire \bridge/conf_pci_am1_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_am1_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[17]/SRNOT ;
    wire \bridge/configuration/pci_addr_mask1[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_am1_out[15]/SRNOT ;
    wire \bridge/conf_pci_am1_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_am1_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[19]/SRNOT ;
    wire \bridge/configuration/pci_addr_mask1[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_addr_mask1[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_am1_out[17]/SRNOT ;
    wire \bridge/conf_pci_am1_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_am1_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFY/SET ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFX/SET ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_sm_bc0_out/SRNOT ;
    wire \bridge/pci_target_unit/pcit_sm_bc0_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/BXNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N360 ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/BXNOT ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N344 ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/BXNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N271 ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFX/SET ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/BXNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N326 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/BYNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_rty_exp_clr/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_conf_offset_out[3]/SRNOT ;
    wire \bridge/pciu_conf_offset_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_conf_offset_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[4]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_conf_offset_out[5]/SRNOT ;
    wire \bridge/pciu_conf_offset_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_conf_offset_out[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_conf_offset_out[7]/SRNOT ;
    wire \bridge/pciu_conf_offset_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pciu_conf_offset_out[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/status_bit8/LOGIC_ONE ;
    wire \bridge/configuration/status_bit8/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[4]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[4]/SRNOT ;
    wire \bridge/configuration/config_addr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[4]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/previous_frame/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/previous_frame/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[6]/SRNOT ;
    wire \bridge/configuration/config_addr[6]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[6]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[7]/SRNOT ;
    wire \bridge/configuration/config_addr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[8]/SRNOT ;
    wire \bridge/configuration/config_addr[8]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_cs_bit31_24[25]/SRNOT ;
    wire \bridge/configuration/pci_err_cs_bit31_24[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_cs_bit31_24[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[10]/SRNOT ;
    wire \bridge/configuration/config_addr[10]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[10]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_cs_bit31_24[27]/SRNOT ;
    wire \bridge/configuration/pci_err_cs_bit31_24[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_cs_bit31_24[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[1]/SRNOT ;
    wire \bridge/configuration/pci_err_data[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[3]/SRNOT ;
    wire \bridge/configuration/pci_err_data[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[5]/SRNOT ;
    wire \bridge/configuration/pci_err_data[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[0]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[0]/BYNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[0]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_waddr[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[7]/SRNOT ;
    wire \bridge/configuration/pci_err_data[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/icr_soft_res/SRNOT ;
    wire \bridge/configuration/icr_soft_res/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[9]/SRNOT ;
    wire \bridge/configuration/pci_err_data[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[1]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[3]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[13]/SRNOT ;
    wire \bridge/configuration/wb_base_addr1[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[21]/SRNOT ;
    wire \bridge/configuration/wb_base_addr1[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[5]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[15]/SRNOT ;
    wire \bridge/configuration/wb_base_addr1[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_ba1_out[19]/SRNOT ;
    wire \bridge/conf_wb_ba1_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_ba1_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[23]/SRNOT ;
    wire \bridge/configuration/wb_base_addr1[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_io_mux/ad_load_ctrl_mhigh/GROM ;
    wire \bridge/pci_io_mux/ad_load_ctrl_mhigh/FROM ;
    wire \bridge/configuration/wb_err_addr[7]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[17]/SRNOT ;
    wire \bridge/configuration/wb_base_addr1[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_ba1_out[13]/SRNOT ;
    wire \bridge/conf_wb_ba1_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_ba1_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[9]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[19]/SRNOT ;
    wire \bridge/configuration/wb_base_addr1[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_base_addr1[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_ba1_out[15]/SRNOT ;
    wire \bridge/conf_wb_ba1_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_ba1_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[13]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[21]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_io_space_enable_out/SRNOT ;
    wire \bridge/conf_io_space_enable_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_ba1_out[17]/SRNOT ;
    wire \bridge/conf_wb_ba1_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_ba1_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[15]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[23]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[31]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_mem_space_enable_out/SRNOT ;
    wire \bridge/conf_mem_space_enable_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_master_enable_out/SRNOT ;
    wire \bridge/conf_pci_master_enable_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[17]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[25]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[19]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[27]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[29]/SRNOT ;
    wire \bridge/configuration/pci_tran_addr1[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_tran_addr1[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_error_en/SRNOT ;
    wire \bridge/configuration/pci_error_en/FFY/ASYNC_FF_GSR_OR ;
    wire \N12330/GROM ;
    wire \bridge/parity_checker/syn3190/GROM ;
    wire \bridge/parity_checker/syn3189/GROM ;
    wire \syn18670/GROM ;
    wire \syn18670/FROM ;
    wire \CRT/ssvga_fifo/gray_read_ptr[1]/SRNOT ;
    wire \CRT/ssvga_fifo/gray_read_ptr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/gray_read_ptr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \syn181997/GROM ;
    wire \syn181997/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[0]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[0]/FROM ;
    wire \CRT/ssvga_fifo/gray_read_ptr[3]/SRNOT ;
    wire \CRT/ssvga_fifo/gray_read_ptr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/gray_read_ptr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \syn182002/GROM ;
    wire \syn182002/FROM ;
    wire \N12313/GROM ;
    wire \N12313/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy/FROM ;
    wire \CRT/ssvga_fifo/gray_read_ptr[5]/SRNOT ;
    wire \CRT/ssvga_fifo/gray_read_ptr[5]/FROM ;
    wire \CRT/ssvga_fifo/gray_read_ptr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/gray_read_ptr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[0]/BYNOT ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[0]/FFY/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/gray_read_ptr[7]/SRNOT ;
    wire \CRT/ssvga_fifo/gray_read_ptr[7]/GROM ;
    wire \CRT/ssvga_fifo/gray_read_ptr[7]/FROM ;
    wire \CRT/ssvga_fifo/gray_read_ptr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/gray_read_ptr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/gray_read_ptr[9]/SRNOT ;
    wire \CRT/ssvga_fifo/gray_read_ptr[9]/FROM ;
    wire \CRT/ssvga_fifo/gray_read_ptr[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/gray_read_ptr[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/BYNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[2]/SRNOT ;
    wire \bridge/configuration/config_addr[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/config_addr[2]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[21]/SRNOT ;
    wire \bridge/configuration/wb_addr_mask1[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[13]/SRNOT ;
    wire \bridge/configuration/wb_addr_mask1[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[23]/SRNOT ;
    wire \bridge/configuration/wb_addr_mask1[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_am1_out[19]/SRNOT ;
    wire \bridge/conf_wb_am1_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_am1_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[15]/SRNOT ;
    wire \bridge/configuration/wb_addr_mask1[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \syn24519/GROM ;
    wire \syn24519/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/req_done_reg/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/req_done_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_am1_out[13]/SRNOT ;
    wire \bridge/conf_wb_am1_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_am1_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[17]/SRNOT ;
    wire \bridge/configuration/wb_addr_mask1[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[19]/SRNOT ;
    wire \bridge/configuration/wb_addr_mask1[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_addr_mask1[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_am1_out[15]/SRNOT ;
    wire \bridge/conf_wb_am1_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_am1_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/delete_wb_err_cs_bit8/SRNOT ;
    wire \bridge/configuration/delete_wb_err_cs_bit8/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/line_end2/SRNOT ;
    wire \CRT/ssvga_crtc/line_end2/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/line_end2/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_am1_out[17]/SRNOT ;
    wire \bridge/conf_wb_am1_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_am1_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[11]/SRNOT ;
    wire \bridge/configuration/wb_err_data[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[21]/SRNOT ;
    wire \bridge/configuration/wb_err_data[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[13]/SRNOT ;
    wire \bridge/configuration/wb_err_data[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[31]/SRNOT ;
    wire \bridge/configuration/wb_err_data[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[23]/SRNOT ;
    wire \bridge/configuration/wb_err_data[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[15]/SRNOT ;
    wire \bridge/configuration/wb_err_data[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[25]/SRNOT ;
    wire \bridge/configuration/wb_err_data[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[17]/SRNOT ;
    wire \bridge/configuration/wb_err_data[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[27]/SRNOT ;
    wire \bridge/configuration/wb_err_data[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[19]/SRNOT ;
    wire \bridge/configuration/wb_err_data[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[29]/SRNOT ;
    wire \bridge/configuration/wb_err_data[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[1]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[3]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[5]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \crt_hsync/BYNOT ;
    wire \crt_hsync/SRNOT ;
    wire \crt_hsync/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[7]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_img_ctrl1_out[0]/SRNOT ;
    wire \bridge/conf_pci_img_ctrl1_out[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[9]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_img_ctrl1[2]/SRNOT ;
    wire \bridge/configuration/pci_img_ctrl1[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_err_pending_out/LOGIC_ONE ;
    wire \bridge/conf_pci_err_pending_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_mem_io1_out/SRNOT ;
    wire \bridge/conf_wb_mem_io1_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_bc_out[2]/LOGIC_ONE ;
    wire \bridge/wishbone_slave_unit/del_sync_bc_out[2]/BXNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_bc_out[2]/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_bc_out[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync_bc_out[2]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_sm_first_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_sm_first_out/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/transfer_input ;
    wire \bridge/wishbone_slave_unit/pcim_sm_first_out/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/CENOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[11]/SRNOT ;
    wire \bridge/configuration/pci_err_data[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/sync_comp_done/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/sync_comp_done/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_done/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_done/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_bc_out[1]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_bc_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_bc_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[21]/SRNOT ;
    wire \bridge/configuration/pci_err_data[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[13]/SRNOT ;
    wire \bridge/configuration/pci_err_data[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_bc_out[3]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_bc_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_bc_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[31]/SRNOT ;
    wire \bridge/configuration/pci_err_data[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[23]/SRNOT ;
    wire \bridge/configuration/pci_err_data[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[15]/SRNOT ;
    wire \bridge/configuration/pci_err_data[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/LOGIC_ONE ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[25]/SRNOT ;
    wire \bridge/configuration/pci_err_data[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[17]/SRNOT ;
    wire \bridge/configuration/pci_err_data[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/LOGIC_ONE ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[27]/SRNOT ;
    wire \bridge/configuration/pci_err_data[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[19]/SRNOT ;
    wire \bridge/configuration/pci_err_data[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/BYNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[29]/SRNOT ;
    wire \bridge/configuration/pci_err_data[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_data[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \N_LED/SRNOT ;
    wire \N_LED/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[11]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[21]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[13]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit31_24[31]/SRNOT ;
    wire \bridge/configuration/wb_err_cs_bit31_24[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit31_24[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[31]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[23]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[15]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit31_24[25]/SRNOT ;
    wire \bridge/configuration/wb_err_cs_bit31_24[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit31_24[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[25]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[17]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit31_24[27]/SRNOT ;
    wire \bridge/configuration/wb_err_cs_bit31_24[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit31_24[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[27]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[19]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/rd_ssvga_en/SRNOT ;
    wire \CRT/ssvga_fifo/rd_ssvga_en/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit31_24[29]/SRNOT ;
    wire \bridge/configuration/wb_err_cs_bit31_24[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_cs_bit31_24[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[29]/SRNOT ;
    wire \bridge/configuration/wb_err_addr[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_addr[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[13]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[21]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_be_out[1]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_be_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_be_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[15]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[31]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[23]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_be_out[3]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_be_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_be_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[17]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[25]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_io_mux/ad_load_ctrl_high/GROM ;
    wire \bridge/pci_io_mux/ad_load_ctrl_high/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[27]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[19]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/sync_req_rty_exp/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/sync_req_rty_exp/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[29]/SRNOT ;
    wire \bridge/configuration/wb_tran_addr1[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_tran_addr1[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/crtc_hblank/SRNOT ;
    wire \CRT/crtc_hblank/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[3]/SRNOT ;
    wire \CRT/pix_start_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[5]/SRNOT ;
    wire \CRT/pix_start_addr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/parity_checker/master_perr_report/SRNOT ;
    wire \bridge/parity_checker/master_perr_report/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_img_ctrl1[2]/SRNOT ;
    wire \bridge/configuration/wb_img_ctrl1[2]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_img_ctrl1[2]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[7]/SRNOT ;
    wire \CRT/pix_start_addr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_img_ctrl1_out[1]/SRNOT ;
    wire \bridge/conf_wb_img_ctrl1_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[9]/SRNOT ;
    wire \CRT/pix_start_addr[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/status_bit15_11[15]/LOGIC_ONE ;
    wire \bridge/configuration/status_bit15_11[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/C6/N18/GROM ;
    wire \CRT/ssvga_fifo/C6/N18/FROM ;
    wire \CRT/ssvga_fifo/C6/N30/GROM ;
    wire \CRT/ssvga_fifo/C6/N30/FROM ;
    wire \CRT/fifo_out[1]/GROM ;
    wire \CRT/fifo_out[1]/FROM ;
    wire \syn176876/GROM ;
    wire \CRT/ssvga_fifo/C6/N42/GROM ;
    wire \CRT/ssvga_fifo/C6/N42/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[11]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/fifo_out[3]/GROM ;
    wire \CRT/fifo_out[3]/FROM ;
    wire \CRT/fifo_out[5]/GROM ;
    wire \CRT/fifo_out[5]/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_sm_rdy_out/SRNOT ;
    wire \bridge/pci_target_unit/pcit_sm_rdy_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[21]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[13]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/fifo_out[7]/GROM ;
    wire \CRT/fifo_out[7]/FROM ;
    wire \bridge/configuration/interrupt_line[1]/SRNOT ;
    wire \bridge/configuration/interrupt_line[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/interrupt_line[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_latency_tim_out[1]/SRNOT ;
    wire \bridge/conf_latency_tim_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_latency_tim_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[31]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[23]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[15]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/interrupt_line[3]/SRNOT ;
    wire \bridge/configuration/interrupt_line[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/interrupt_line[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_latency_tim_out[3]/SRNOT ;
    wire \bridge/conf_latency_tim_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_latency_tim_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[25]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[17]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/interrupt_line[5]/SRNOT ;
    wire \bridge/configuration/interrupt_line[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/interrupt_line[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_latency_tim_out[5]/SRNOT ;
    wire \bridge/conf_latency_tim_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_latency_tim_out[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[27]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[19]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/BYNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/interrupt_line[7]/SRNOT ;
    wire \bridge/configuration/interrupt_line[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/interrupt_line[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/int_prop_en/SRNOT ;
    wire \bridge/configuration/int_prop_en/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_latency_tim_out[7]/SRNOT ;
    wire \bridge/conf_latency_tim_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_latency_tim_out[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/error_int_en/SRNOT ;
    wire \bridge/configuration/error_int_en/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[29]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/perr_int_en/SRNOT ;
    wire \bridge/configuration/perr_int_en/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[21]/SRNOT ;
    wire \bridge/configuration/pci_base_addr1[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[13]/SRNOT ;
    wire \bridge/configuration/pci_base_addr1[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/serr_int_en/SRNOT ;
    wire \bridge/configuration/serr_int_en/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba1_out[19]/SRNOT ;
    wire \bridge/conf_pci_ba1_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba1_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[23]/SRNOT ;
    wire \bridge/configuration/pci_base_addr1[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[15]/SRNOT ;
    wire \bridge/configuration/pci_base_addr1[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba1_out[13]/SRNOT ;
    wire \bridge/conf_pci_ba1_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba1_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[17]/SRNOT ;
    wire \bridge/configuration/pci_base_addr1[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[1]/SRNOT ;
    wire \bridge/configuration/wb_err_data[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy/FROM ;
    wire \bridge/conf_pci_ba1_out[15]/SRNOT ;
    wire \bridge/conf_pci_ba1_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba1_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[19]/SRNOT ;
    wire \bridge/configuration/pci_base_addr1[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr1[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[3]/SRNOT ;
    wire \bridge/configuration/wb_err_data[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba1_out[17]/SRNOT ;
    wire \bridge/conf_pci_ba1_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba1_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[5]/SRNOT ;
    wire \bridge/configuration/wb_err_data[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[7]/SRNOT ;
    wire \bridge/configuration/wb_err_data[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \syn22225/GROM ;
    wire \syn22225/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[9]/SRNOT ;
    wire \bridge/configuration/wb_err_data[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/wb_err_data[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \syn181402/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/GROM ;
    wire N12592;
    wire \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wbu_mabort_rec_out/SRNOT ;
    wire \bridge/wbu_mabort_rec_out/GROM ;
    wire \bridge/wbu_mabort_rec_out/FROM ;
    wire \bridge/wbu_mabort_rec_out/FFX/ASYNC_FF_GSR_OR ;
    wire \N12380/GROM ;
    wire \N12380/FROM ;
    wire \N12607/GROM ;
    wire \N12607/FROM ;
    wire \syn18930/GROM ;
    wire \syn18930/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/GROM ;
    wire N12593;
    wire \bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[4]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \syn181005/GROM ;
    wire \syn181005/FROM ;
    wire \N12466/GROM ;
    wire \N12466/FROM ;
    wire \syn181040/GROM ;
    wire \syn181040/FROM ;
    wire \syn178588/GROM ;
    wire \syn178588/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[14]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[14]/FROM ;
    wire \syn181092/GROM ;
    wire \syn181092/FROM ;
    wire \syn181039/GROM ;
    wire \syn181039/FROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[0]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[0]/FROM ;
    wire \CRT/ssvga_wbm_if/N1531/GROM ;
    wire N12635;
    wire \CRT/ssvga_wbm_if/N1531/XORF ;
    wire \syn181347/GROM ;
    wire \syn17084/GROM ;
    wire \syn17084/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[0]/GROM ;
    wire \syn179378/GROM ;
    wire \syn180806/GROM ;
    wire \syn180806/FROM ;
    wire \syn181107/GROM ;
    wire \syn181107/FROM ;
    wire \syn19708/GROM ;
    wire \syn19562/GROM ;
    wire \syn19562/FROM ;
    wire \syn179377/GROM ;
    wire \syn60043/GROM ;
    wire \syn60043/FROM ;
    wire \syn60048/GROM ;
    wire \syn60048/FROM ;
    wire \syn17119/GROM ;
    wire \syn17119/FROM ;
    wire \rgb_int[10]/GROM ;
    wire \rgb_int[10]/FROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C707/GROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/C707/FROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[2]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[2]/FROM ;
    wire \syn180469/GROM ;
    wire \syn180469/FROM ;
    wire \syn16983/GROM ;
    wire \syn16983/FROM ;
    wire \syn60047/GROM ;
    wire \syn60047/FROM ;
    wire \syn181605/GROM ;
    wire \syn181605/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/ad_en_w/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/ad_en_w/FROM ;
    wire \CRT/ssvga_fifo/S_43/cell0/GROM ;
    wire \rgb_int[8]/GROM ;
    wire \rgb_int[8]/FROM ;
    wire \syn180794/GROM ;
    wire \syn180794/FROM ;
    wire \syn17017/GROM ;
    wire \syn17017/FROM ;
    wire \syn182602/GROM ;
    wire \syn182602/FROM ;
    wire \syn180467/GROM ;
    wire \syn180467/FROM ;
    wire \syn180843/GROM ;
    wire \syn180843/FROM ;
    wire \syn180939/GROM ;
    wire \syn180939/FROM ;
    wire \syn182601/GROM ;
    wire \syn182601/FROM ;
    wire \rgb_int[6]/GROM ;
    wire \rgb_int[6]/FROM ;
    wire \rgb_int[14]/GROM ;
    wire \rgb_int[14]/FROM ;
    wire \syn20874/GROM ;
    wire \syn180466/GROM ;
    wire \syn180466/FROM ;
    wire \syn180658/GROM ;
    wire \syn180658/FROM ;
    wire \syn180763/GROM ;
    wire \syn180763/FROM ;
    wire \syn180792/GROM ;
    wire \syn180792/FROM ;
    wire \syn180938/GROM ;
    wire \syn180938/FROM ;
    wire \syn181145/GROM ;
    wire \syn181145/FROM ;
    wire \syn182473/GROM ;
    wire \syn182473/FROM ;
    wire \syn182628/GROM ;
    wire \syn182663/GROM ;
    wire \syn182663/FROM ;
    wire \syn178884/GROM ;
    wire \syn178884/FROM ;
    wire \bridge/pci_target_unit/pci_target_if/n_1317/GROM ;
    wire \bridge/pci_target_unit/pci_target_if/n_1317/FROM ;
    wire \syn180657/GROM ;
    wire \syn180657/FROM ;
    wire \syn180937/GROM ;
    wire \syn180937/FROM ;
    wire \syn181144/GROM ;
    wire \syn181144/FROM ;
    wire \syn20872/GROM ;
    wire \syn20872/FROM ;
    wire \syn182627/GROM ;
    wire \syn182662/GROM ;
    wire \syn182662/FROM ;
    wire \bridge/pci_target_unit/fifos/pciw_rallow/GROM ;
    wire \bridge/pci_target_unit/fifos/pciw_rallow/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[16]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[16]/FROM ;
    wire \syn17052/GROM ;
    wire \syn17052/FROM ;
    wire \rgb_int[4]/GROM ;
    wire \rgb_int[4]/FROM ;
    wire \rgb_int[12]/GROM ;
    wire \rgb_int[12]/FROM ;
    wire \syn180523/GROM ;
    wire \syn180523/FROM ;
    wire \syn180841/GROM ;
    wire \syn180841/FROM ;
    wire \syn180957/GROM ;
    wire \syn180957/FROM ;
    wire \syn179985/GROM ;
    wire \syn179985/FROM ;
    wire \syn120400/GROM ;
    wire \syn120400/FROM ;
    wire \N12478/GROM ;
    wire \N12478/FROM ;
    wire \syn182610/GROM ;
    wire \syn182610/FROM ;
    wire \syn177733/GROM ;
    wire \syn177733/FROM ;
    wire \syn16919/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[17]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[17]/FROM ;
    wire \syn180522/GROM ;
    wire \syn180522/FROM ;
    wire \syn180701/GROM ;
    wire \syn180701/FROM ;
    wire \syn21246/GROM ;
    wire \syn21246/FROM ;
    wire \syn180669/GROM ;
    wire \syn180669/FROM ;
    wire \bridge/configuration/C287/N3/GROM ;
    wire \bridge/configuration/C287/N3/FROM ;
    wire \syn18659/GROM ;
    wire \syn18659/FROM ;
    wire \syn16939/GROM ;
    wire \syn16939/FROM ;
    wire \syn17875/GROM ;
    wire \syn17875/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[26]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[26]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[18]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[18]/FROM ;
    wire \syn180521/GROM ;
    wire \syn180521/FROM ;
    wire \syn180700/GROM ;
    wire \syn180700/FROM ;
    wire \syn180840/GROM ;
    wire \syn180840/FROM ;
    wire \syn180951/GROM ;
    wire \syn180951/FROM ;
    wire \syn17971/GROM ;
    wire \syn17971/FROM ;
    wire \syn181166/GROM ;
    wire \syn181166/FROM ;
    wire \syn177524/GROM ;
    wire \syn177524/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en/GROM ;
    wire \syn177830/GROM ;
    wire \syn177830/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[28]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[28]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[27]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[27]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[19]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[19]/FROM ;
    wire \syn180699/GROM ;
    wire \syn180699/FROM ;
    wire \syn181194/GROM ;
    wire \syn181194/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/cnf_progress/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/cnf_progress/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/cnf_progress/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/cnf_progress/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[22]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[22]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[4]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[4]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[28]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[28]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[20]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[20]/FROM ;
    wire \syn180205/GROM ;
    wire \syn180205/FROM ;
    wire \syn180660/GROM ;
    wire \syn180660/FROM ;
    wire \syn21571/GROM ;
    wire \syn21571/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[12]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[12]/FROM ;
    wire \syn178999/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[6]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[6]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[29]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[29]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[21]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[21]/FROM ;
    wire \syn179931/GROM ;
    wire \syn179931/FROM ;
    wire \syn180138/GROM ;
    wire \syn180138/FROM ;
    wire \syn20484/GROM ;
    wire \syn20484/FROM ;
    wire \syn178054/GROM ;
    wire \syn178054/FROM ;
    wire \syn180884/GROM ;
    wire \syn180884/FROM ;
    wire \syn180907/GROM ;
    wire \syn180907/FROM ;
    wire \syn181146/GROM ;
    wire \syn181146/FROM ;
    wire \syn181403/GROM ;
    wire \syn182474/GROM ;
    wire \syn182474/FROM ;
    wire \syn17073/GROM ;
    wire \syn17073/FROM ;
    wire \syn18756/GROM ;
    wire \syn178848/GROM ;
    wire \syn178848/FROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[24]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[24]/FROM ;
    wire \syn178998/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[30]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[30]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[22]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[22]/FROM ;
    wire \syn178236/GROM ;
    wire \syn178236/FROM ;
    wire \syn20909/GROM ;
    wire \syn20909/FROM ;
    wire \syn20934/GROM ;
    wire \syn20934/FROM ;
    wire \syn177954/GROM ;
    wire \syn177954/FROM ;
    wire \syn180626/GROM ;
    wire \syn180626/FROM ;
    wire \syn177921/GROM ;
    wire \syn177921/FROM ;
    wire \syn179848/GROM ;
    wire \syn179848/FROM ;
    wire \N12311/GROM ;
    wire \N12311/FROM ;
    wire \syn182394/GROM ;
    wire \syn182394/FROM ;
    wire \syn182432/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[16]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[16]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[7]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[7]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[31]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[31]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[23]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[23]/FROM ;
    wire \syn180122/GROM ;
    wire \syn180122/FROM ;
    wire \syn120384/GROM ;
    wire \syn178092/GROM ;
    wire \syn178092/FROM ;
    wire \syn120382/GROM ;
    wire \syn120382/FROM ;
    wire \syn20770/GROM ;
    wire \syn20770/FROM ;
    wire \syn182423/GROM ;
    wire \syn182423/FROM ;
    wire \syn178179/GROM ;
    wire \syn178179/FROM ;
    wire \syn24474/GROM ;
    wire \syn24474/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[25]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[25]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[17]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[17]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[8]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[8]/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/S_291/cell0/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/S_291/cell0/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[24]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[24]/FROM ;
    wire \syn16934/GROM ;
    wire \syn16934/FROM ;
    wire \syn180098/GROM ;
    wire \syn180098/FROM ;
    wire \syn180121/GROM ;
    wire \syn180121/FROM ;
    wire \syn21091/GROM ;
    wire \syn21091/FROM ;
    wire \syn60044/GROM ;
    wire \syn60044/FROM ;
    wire \syn18468/GROM ;
    wire \syn18468/FROM ;
    wire \syn17071/GROM ;
    wire \syn17071/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[26]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[26]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[18]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[18]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[9]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[9]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[1]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[1]/FROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[25]/GROM ;
    wire \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[25]/FROM ;
    wire \syn17102/GROM ;
    wire \syn17102/FROM ;
    wire \syn20773/GROM ;
    wire \syn20773/FROM ;
    wire \syn180420/GROM ;
    wire \syn180420/FROM ;
    wire \syn181037/GROM ;
    wire \syn181037/FROM ;
    wire \syn182526/GROM ;
    wire \syn178201/GROM ;
    wire \syn178201/FROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[28]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[28]/FROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[20]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[20]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[10]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[10]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[2]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[2]/FROM ;
    wire \syn178436/GROM ;
    wire \syn178436/FROM ;
    wire \syn179850/GROM ;
    wire \syn179850/FROM ;
    wire \syn21507/GROM ;
    wire \syn21507/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/C983/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/C983/FROM ;
    wire \syn182535/GROM ;
    wire \syn182535/FROM ;
    wire \syn182555/GROM ;
    wire \syn182555/FROM ;
    wire \syn18965/GROM ;
    wire \syn18965/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[22]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[22]/FROM ;
    wire \bridge/pci_target_unit/fifos/out_count_en/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[12]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[12]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[3]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[3]/FROM ;
    wire \bridge/configuration/C292/N3/GROM ;
    wire \bridge/configuration/C292/N3/FROM ;
    wire \syn179878/GROM ;
    wire \syn179878/FROM ;
    wire \syn20740/GROM ;
    wire \syn20740/FROM ;
    wire \syn179950/GROM ;
    wire \syn179950/FROM ;
    wire \syn20769/GROM ;
    wire \syn20769/FROM ;
    wire \syn180611/GROM ;
    wire \syn180611/FROM ;
    wire \syn177820/GROM ;
    wire \syn177820/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/load_force/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/load_force/FROM ;
    wire \syn18944/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[30]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[30]/FROM ;
    wire \bridge/pci_target_unit/pci_target_if/n_1298/GROM ;
    wire \bridge/pci_target_unit/pci_target_if/n_1298/FROM ;
    wire \bridge/configuration/C346/N5/GROM ;
    wire \bridge/configuration/C346/N5/FROM ;
    wire \bridge/configuration/C284/N39/GROM ;
    wire \bridge/configuration/C284/N39/FROM ;
    wire \syn179912/GROM ;
    wire \syn179912/FROM ;
    wire \syn178200/GROM ;
    wire \syn178200/FROM ;
    wire \syn120386/GROM ;
    wire \syn120386/FROM ;
    wire \bridge/pci_target_unit/pci_target_if/n_1335/GROM ;
    wire \bridge/pci_target_unit/pci_target_if/n_1335/FROM ;
    wire \syn18655/GROM ;
    wire \syn18655/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[13]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[13]/FROM ;
    wire \syn178433/GROM ;
    wire \syn178433/FROM ;
    wire \syn180107/GROM ;
    wire \syn180107/FROM ;
    wire \syn180609/GROM ;
    wire \syn180609/FROM ;
    wire \syn17031/GROM ;
    wire \syn17031/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[5]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[5]/FROM ;
    wire \syn17023/GROM ;
    wire \syn17023/FROM ;
    wire \bridge/pci_target_unit/del_sync/comp_rty_exp_reg/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/comp_rty_exp_reg/GROM ;
    wire N12602;
    wire \bridge/pci_target_unit/del_sync/comp_rty_exp_reg/FFX/ASYNC_FF_GSR_OR ;
    wire \syn17895/GROM ;
    wire \syn17895/FROM ;
    wire \syn178106/GROM ;
    wire \syn178106/FROM ;
    wire \syn178356/GROM ;
    wire \syn178356/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N40 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow/FROM ;
    wire \syn17005/GROM ;
    wire \bridge/configuration/C285/N99/GROM ;
    wire \bridge/configuration/C285/N99/FROM ;
    wire \bridge/configuration/C296/N24/GROM ;
    wire \bridge/configuration/C296/N24/FROM ;
    wire \bridge/configuration/C293/N14/GROM ;
    wire \bridge/configuration/C293/N14/FROM ;
    wire \syn180261/GROM ;
    wire \syn180261/FROM ;
    wire \bridge/configuration/C286/N19/GROM ;
    wire \bridge/configuration/C286/N19/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[21]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[21]/FROM ;
    wire \syn182037/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/read_completed_reg/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_sm/read_completed_reg/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/read_completed_reg/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/read_completed_reg/FFX/ASYNC_FF_GSR_OR ;
    wire \syn177990/GROM ;
    wire \syn177990/FROM ;
    wire \syn24470/GROM ;
    wire \syn24470/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[24]/GROM ;
    wire \bridge/configuration/C298/N3/GROM ;
    wire \bridge/configuration/C298/N3/FROM ;
    wire \syn179762/GROM ;
    wire \syn179762/FROM ;
    wire \syn178462/GROM ;
    wire \syn178462/FROM ;
    wire \syn178883/GROM ;
    wire \syn178883/FROM ;
    wire \syn180316/GROM ;
    wire \syn180316/FROM ;
    wire \syn17120/GROM ;
    wire \syn17120/FROM ;
    wire \syn180270/GROM ;
    wire \syn180270/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[23]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[23]/FROM ;
    wire \N12541/GROM ;
    wire \N12541/FROM ;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_reg/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_reg/FROM ;
    wire \bridge/pci_target_unit/del_sync/req_rty_exp_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \syn177989/GROM ;
    wire \syn177989/FROM ;
    wire \syn177710/GROM ;
    wire \syn177710/FROM ;
    wire \bridge/configuration/C294/N29/GROM ;
    wire \bridge/configuration/C294/N29/FROM ;
    wire \syn180315/GROM ;
    wire \syn180315/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[11]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[11]/FROM ;
    wire \syn177922/GROM ;
    wire \syn177922/FROM ;
    wire \syn178094/GROM ;
    wire \syn178094/FROM ;
    wire \syn178311/GROM ;
    wire \syn178311/FROM ;
    wire \syn179789/GROM ;
    wire \syn180314/GROM ;
    wire \syn180314/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[27]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[27]/FROM ;
    wire \syn17077/GROM ;
    wire \syn17077/FROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[3]/GROM ;
    wire \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[3]/FROM ;
    wire \bridge/configuration/C290/N99/GROM ;
    wire \bridge/configuration/C290/N99/FROM ;
    wire \syn21466/GROM ;
    wire \syn21466/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[15]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[15]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[29]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[29]/FROM ;
    wire \syn17056/GROM ;
    wire \syn177925/GROM ;
    wire \syn177925/FROM ;
    wire \syn177869/GROM ;
    wire \syn177869/FROM ;
    wire \syn18087/GROM ;
    wire \syn18087/FROM ;
    wire \syn24466/GROM ;
    wire \syn24466/FROM ;
    wire \syn16984/GROM ;
    wire \syn16984/FROM ;
    wire \syn178535/GROM ;
    wire \syn178535/FROM ;
    wire \bridge/configuration/C296/N64/GROM ;
    wire \bridge/configuration/C296/N64/FROM ;
    wire \bridge/configuration/C297/N84/GROM ;
    wire \bridge/configuration/C297/N84/FROM ;
    wire \syn179761/GROM ;
    wire \syn179761/FROM ;
    wire \syn179847/GROM ;
    wire \syn179847/FROM ;
    wire \syn179894/GROM ;
    wire \syn180052/GROM ;
    wire \syn180052/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[30]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[30]/FROM ;
    wire \syn17020/GROM ;
    wire \syn17020/FROM ;
    wire \syn178035/GROM ;
    wire \syn178035/FROM ;
    wire \syn178240/GROM ;
    wire \syn178240/FROM ;
    wire \syn19064/GROM ;
    wire \syn19064/FROM ;
    wire \bridge/configuration/C291/N14/GROM ;
    wire \bridge/configuration/C291/N14/FROM ;
    wire \syn18784/GROM ;
    wire \syn18784/FROM ;
    wire \syn179948/GROM ;
    wire \syn179948/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/C103/N15 ;
    wire \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/FFX/ASYNC_FF_GSR_OR ;
    wire \syn177613/GROM ;
    wire \syn177613/FROM ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy/GROM ;
    wire \bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy/FROM ;
    wire \syn178376/GROM ;
    wire \syn178376/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[19]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_sm_data_out[19]/FROM ;
    wire \syn178132/GROM ;
    wire \syn178132/FROM ;
    wire \syn18717/GROM ;
    wire \syn18717/FROM ;
    wire \bridge/configuration/C294/N84/GROM ;
    wire \bridge/configuration/C294/N84/FROM ;
    wire \bridge/configuration/C294/N69/GROM ;
    wire \bridge/configuration/C294/N69/FROM ;
    wire \bridge/configuration/C297/N69/GROM ;
    wire \bridge/configuration/C297/N69/FROM ;
    wire \bridge/pci_target_unit/del_sync/comp_done_reg_clr/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/comp_done_reg_clr/FFY/ASYNC_FF_GSR_OR ;
    wire \syn177655/GROM ;
    wire \syn177655/FROM ;
    wire \syn177670/GROM ;
    wire \syn177670/FROM ;
    wire \syn178058/GROM ;
    wire \syn178058/FROM ;
    wire \syn178131/GROM ;
    wire \syn178131/FROM ;
    wire \syn18567/GROM ;
    wire \syn18567/FROM ;
    wire \syn177732/GROM ;
    wire \syn177732/FROM ;
    wire \syn18681/GROM ;
    wire \syn18681/FROM ;
    wire \syn20277/GROM ;
    wire \syn20277/FROM ;
    wire \bridge/configuration/C286/N54/GROM ;
    wire \bridge/configuration/C286/N54/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C262/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C262/FROM ;
    wire \syn178394/GROM ;
    wire \syn178394/FROM ;
    wire \syn59929/GROM ;
    wire \syn59929/FROM ;
    wire \syn178313/GROM ;
    wire \syn178514/GROM ;
    wire \syn179544/GROM ;
    wire \syn19914/GROM ;
    wire \syn19914/FROM ;
    wire \syn17080/GROM ;
    wire \syn17080/FROM ;
    wire \syn16988/GROM ;
    wire \N12163/GROM ;
    wire \N12163/FROM ;
    wire \N12152/GROM ;
    wire \syn20367/GROM ;
    wire \syn20367/FROM ;
    wire \N12312/GROM ;
    wire \N12312/FROM ;
    wire \syn17054/GROM ;
    wire \syn177790/GROM ;
    wire \syn177790/FROM ;
    wire \bridge/configuration/C286/N99/GROM ;
    wire \bridge/configuration/C286/N99/FROM ;
    wire \syn17856/GROM ;
    wire \syn17856/FROM ;
    wire \syn177693/GROM ;
    wire \syn177693/FROM ;
    wire \syn177857/GROM ;
    wire \syn177857/FROM ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/C0/C116/GROM ;
    wire \syn177574/GROM ;
    wire \syn177574/FROM ;
    wire \syn18010/GROM ;
    wire \syn18010/FROM ;
    wire \syn177856/GROM ;
    wire \syn177856/FROM ;
    wire \syn60060/GROM ;
    wire \syn60060/FROM ;
    wire \syn177609/GROM ;
    wire \syn177609/FROM ;
    wire \syn178055/GROM ;
    wire \syn178055/FROM ;
    wire \syn48756/GROM ;
    wire \syn50321/GROM ;
    wire \syn177657/GROM ;
    wire \syn177657/FROM ;
    wire \syn177778/GROM ;
    wire \syn177778/FROM ;
    wire \syn17990/GROM ;
    wire \syn17990/FROM ;
    wire \syn60089/GROM ;
    wire \syn60089/FROM ;
    wire \syn60045/GROM ;
    wire \syn60045/FROM ;
    wire \syn177568/GROM ;
    wire \syn177585/GROM ;
    wire \syn177585/FROM ;
    wire \syn177738/GROM ;
    wire \syn177738/FROM ;
    wire \syn17057/GROM ;
    wire \N12065/GROM ;
    wire \N12065/FROM ;
    wire \syn17004/GROM ;
    wire \syn17004/FROM ;
    wire \syn177501/GROM ;
    wire \syn177501/FROM ;
    wire \syn177608/GROM ;
    wire \syn177608/FROM ;
    wire \syn177569/GROM ;
    wire \syn177656/GROM ;
    wire \syn177656/FROM ;
    wire \syn17115/GROM ;
    wire \syn17115/FROM ;
    wire \bridge/configuration/wb_error_en/SRNOT ;
    wire \bridge/configuration/wb_error_en/FFY/ASYNC_FF_GSR_OR ;
    wire \syn177260/GROM ;
    wire \syn177260/FROM ;
    wire \syn177541/GROM ;
    wire \syn18051/GROM ;
    wire \CRT/ssvga_fifo/C6/N6/GROM ;
    wire \CRT/ssvga_fifo/C6/N6/FROM ;
    wire \syn176894/GROM ;
    wire \syn176894/FROM ;
    wire \syn177406/GROM ;
    wire \syn177406/FROM ;
    wire \syn177563/GROM ;
    wire \syn177563/FROM ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/C0/C112/GROM ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/C0/C112/FROM ;
    wire \bridge/pci_mux_par_in/GROM ;
    wire \bridge/configuration/pci_base_addr0[21]/SRNOT ;
    wire \bridge/configuration/pci_base_addr0[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[13]/SRNOT ;
    wire \bridge/configuration/pci_base_addr0[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/sync_req_comp_pending/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/sync_req_comp_pending/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba0_out[19]/SRNOT ;
    wire \bridge/conf_pci_ba0_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba0_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[23]/SRNOT ;
    wire \bridge/configuration/pci_base_addr0[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[15]/SRNOT ;
    wire \bridge/configuration/pci_base_addr0[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_wb_err_pending_out/LOGIC_ONE ;
    wire \bridge/conf_wb_err_pending_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba0_out[13]/SRNOT ;
    wire \bridge/conf_pci_ba0_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba0_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[17]/SRNOT ;
    wire \bridge/configuration/pci_base_addr0[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[19]/SRNOT ;
    wire \bridge/configuration/pci_base_addr0[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_base_addr0[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba0_out[15]/SRNOT ;
    wire \bridge/conf_pci_ba0_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba0_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba0_out[17]/SRNOT ;
    wire \bridge/conf_pci_ba0_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_ba0_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/BYNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[1]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[3]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[5]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/status_bit15_11[14]/LOGIC_ONE ;
    wire \bridge/configuration/status_bit15_11[14]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[7]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[9]/SRNOT ;
    wire \bridge/configuration/pci_err_addr[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/pci_err_addr[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/status_bit15_11[13]/LOGIC_ONE ;
    wire \bridge/configuration/status_bit15_11[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/configuration/status_bit15_11[12]/LOGIC_ONE ;
    wire \bridge/configuration/status_bit15_11[12]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[11]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFY/SET ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[21]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[13]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFX/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[31]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[23]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[15]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFY/RST ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFX/SET ;
    wire \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[25]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[17]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_pci_mem_io1_out/SRNOT ;
    wire \bridge/conf_pci_mem_io1_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/parity_checker/BLK0_4/GROM ;
    wire \bridge/parity_checker/syn3234 ;
    wire \bridge/parity_checker/BLK0_4/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[11]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/parity_checker/BLK1_4/CYINIT ;
    wire \bridge/parity_checker/BLK1_4/GROM ;
    wire \bridge/parity_checker/syn3232 ;
    wire \bridge/parity_checker/BLK1_4/XORF ;
    wire \bridge/parity_checker/BLK2_4/CYINIT ;
    wire \bridge/parity_checker/BLK2_4/GROM ;
    wire \bridge/parity_checker/syn3230 ;
    wire \bridge/parity_checker/BLK2_4/XORF ;
    wire \bridge/configuration/status_bit15_11[11]/LOGIC_ONE ;
    wire \bridge/configuration/status_bit15_11[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/parity_checker/BLK3_4/GROM ;
    wire \bridge/parity_checker/syn3228 ;
    wire \bridge/parity_checker/BLK3_4/XORF ;
    wire \bridge/parity_checker/BLK4_4/CYINIT ;
    wire \bridge/parity_checker/BLK4_4/GROM ;
    wire \bridge/parity_checker/syn3226 ;
    wire \bridge/parity_checker/BLK4_4/XORF ;
    wire \CRT/pix_start_addr[11]/SRNOT ;
    wire \CRT/pix_start_addr[11]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[11]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/parity_checker/par_gen/syn156 ;
    wire \bridge/parity_checker/par_gen/BLK0_2/XORF ;
    wire \RST/IBUF ;
    wire \RST/KEEPER ;
    wire \AD[27]/SRNOT ;
    wire \AD[27]/IDELAY ;
    wire \AD[27]/OD ;
    wire \AD[27]/ENABLE ;
    wire \AD[27]/KEEPER ;
    wire \AD[27]/OUTBUF_GTS_AND ;
    wire \AD[27]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[27]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[27]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[26]/SRNOT ;
    wire \AD[26]/IDELAY ;
    wire \AD[26]/OD ;
    wire \AD[26]/ENABLE ;
    wire \AD[26]/KEEPER ;
    wire \AD[26]/OUTBUF_GTS_AND ;
    wire \AD[26]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[26]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[26]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[25]/SRNOT ;
    wire \AD[25]/IDELAY ;
    wire \AD[25]/OD ;
    wire \AD[25]/ENABLE ;
    wire \AD[25]/KEEPER ;
    wire \AD[25]/OUTBUF_GTS_AND ;
    wire \AD[25]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[25]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[25]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[24]/SRNOT ;
    wire \AD[24]/IDELAY ;
    wire \AD[24]/OD ;
    wire \AD[24]/ENABLE ;
    wire \AD[24]/KEEPER ;
    wire \AD[24]/OUTBUF_GTS_AND ;
    wire \AD[24]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[24]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[24]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[23]/SRNOT ;
    wire \AD[23]/IDELAY ;
    wire \AD[23]/OD ;
    wire \AD[23]/ENABLE ;
    wire \AD[23]/KEEPER ;
    wire \AD[23]/OUTBUF_GTS_AND ;
    wire \AD[23]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[23]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[23]/TFF/ASYNC_FF_GSR_OR ;
    wire \CBE[3]/SRNOT ;
    wire \CBE[3]/IBUF ;
    wire \CBE[3]/IDELAY ;
    wire \CBE[3]/OD ;
    wire \CBE[3]/TNOT ;
    wire \CBE[3]/ENABLE ;
    wire \CBE[3]/KEEPER ;
    wire \CBE[3]/OUTBUF_GTS_AND ;
    wire \CBE[3]/IFF/ASYNC_FF_GSR_OR ;
    wire \CBE[3]/OFF/ASYNC_FF_GSR_OR ;
    wire \CBE[3]/TFF/ASYNC_FF_GSR_OR ;
    wire \IDSEL/IBUF ;
    wire \IDSEL/KEEPER ;
    wire \AD[17]/SRNOT ;
    wire \AD[17]/IDELAY ;
    wire \AD[17]/ENABLE ;
    wire \AD[17]/KEEPER ;
    wire \AD[17]/OUTBUF_GTS_AND ;
    wire \AD[17]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[17]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[17]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[16]/SRNOT ;
    wire \AD[16]/IDELAY ;
    wire \AD[16]/OD ;
    wire \AD[16]/ENABLE ;
    wire \AD[16]/KEEPER ;
    wire \AD[16]/OUTBUF_GTS_AND ;
    wire \AD[16]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[16]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[16]/TFF/ASYNC_FF_GSR_OR ;
    wire \CBE[2]/SRNOT ;
    wire \CBE[2]/IBUF ;
    wire \CBE[2]/IDELAY ;
    wire \CBE[2]/OD ;
    wire \CBE[2]/TNOT ;
    wire \CBE[2]/ENABLE ;
    wire \CBE[2]/KEEPER ;
    wire \CBE[2]/OUTBUF_GTS_AND ;
    wire \CBE[2]/IFF/ASYNC_FF_GSR_OR ;
    wire \CBE[2]/OFF/ASYNC_FF_GSR_OR ;
    wire \CBE[2]/TFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[27]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \STOP/SRNOT ;
    wire \STOP/IBUF ;
    wire \STOP/IDELAY ;
    wire STOP_out;
    wire \STOP/TNOT ;
    wire STOP_en;
    wire \STOP/ENABLE ;
    wire \STOP/KEEPER ;
    wire \STOP/OUTBUF_GTS_AND ;
    wire \STOP/IFF/ASYNC_FF_GSR_OR ;
    wire \STOP/OFF/ASYNC_FF_GSR_OR ;
    wire \STOP/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[22]/SRNOT ;
    wire \AD[22]/IDELAY ;
    wire \AD[22]/OD ;
    wire \AD[22]/ENABLE ;
    wire \AD[22]/KEEPER ;
    wire \AD[22]/OUTBUF_GTS_AND ;
    wire \AD[22]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[22]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[22]/TFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[19]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \FRAME/SRNOT ;
    wire \FRAME/IBUF ;
    wire \FRAME/IDELAY ;
    wire FRAME_out;
    wire \FRAME/TNOT ;
    wire FRAME_en;
    wire \FRAME/ENABLE ;
    wire \FRAME/KEEPER ;
    wire \FRAME/OUTBUF_GTS_AND ;
    wire \FRAME/IFF/ASYNC_FF_GSR_OR ;
    wire \FRAME/OFF/ASYNC_FF_GSR_OR ;
    wire \FRAME/TFF/ASYNC_FF_GSR_OR ;
    wire \PERR/SRNOT ;
    wire \PERR/IBUF ;
    wire \PERR/OD ;
    wire PERR_out;
    wire PERR_en;
    wire \PERR/ENABLE ;
    wire \PERR/KEEPER ;
    wire \PERR/OUTBUF_GTS_AND ;
    wire \PERR/OFF/ASYNC_FF_GSR_OR ;
    wire \PERR/TFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[21]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \AD[21]/SRNOT ;
    wire \AD[21]/IDELAY ;
    wire \AD[21]/OD ;
    wire \AD[21]/ENABLE ;
    wire \AD[21]/KEEPER ;
    wire \AD[21]/OUTBUF_GTS_AND ;
    wire \AD[21]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[21]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[21]/TFF/ASYNC_FF_GSR_OR ;
    wire \IRDY/SRNOT ;
    wire \IRDY/IBUF ;
    wire \IRDY/IDELAY ;
    wire IRDY_out;
    wire \IRDY/TNOT ;
    wire IRDY_en;
    wire \IRDY/ENABLE ;
    wire \IRDY/KEEPER ;
    wire \IRDY/OUTBUF_GTS_AND ;
    wire \IRDY/IFF/ASYNC_FF_GSR_OR ;
    wire \IRDY/OFF/ASYNC_FF_GSR_OR ;
    wire \IRDY/TFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[13]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \AD[20]/SRNOT ;
    wire \AD[20]/IDELAY ;
    wire \AD[20]/OD ;
    wire \AD[20]/ENABLE ;
    wire \AD[20]/KEEPER ;
    wire \AD[20]/OUTBUF_GTS_AND ;
    wire \AD[20]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[20]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[20]/TFF/ASYNC_FF_GSR_OR ;
    wire \SERR/SRNOT ;
    wire \SERR/OD ;
    wire SERR_out;
    wire \SERR/TNOT ;
    wire SERR_en;
    wire \SERR/ENABLE ;
    wire \SERR/KEEPER ;
    wire \SERR/OUTBUF_GTS_AND ;
    wire \SERR/OFF/ASYNC_FF_GSR_OR ;
    wire \SERR/TFF/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[21]/SRNOT ;
    wire \CRT/pix_start_addr[21]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[21]/FFX/ASYNC_FF_GSR_OR ;
    wire \AD[19]/SRNOT ;
    wire \AD[19]/IDELAY ;
    wire \AD[19]/OD ;
    wire \AD[19]/ENABLE ;
    wire \AD[19]/KEEPER ;
    wire \AD[19]/OUTBUF_GTS_AND ;
    wire \AD[19]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[19]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[19]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[13]/SRNOT ;
    wire \AD[13]/IDELAY ;
    wire \AD[13]/OD ;
    wire \AD[13]/ENABLE ;
    wire \AD[13]/KEEPER ;
    wire \AD[13]/OUTBUF_GTS_AND ;
    wire \AD[13]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[13]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[13]/TFF/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[13]/SRNOT ;
    wire \CRT/pix_start_addr[13]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[13]/FFX/ASYNC_FF_GSR_OR ;
    wire \PAR/SRNOT ;
    wire \PAR/IBUF ;
    wire PAR_out;
    wire \PAR/TNOT ;
    wire PAR_en;
    wire \PAR/ENABLE ;
    wire \PAR/KEEPER ;
    wire \PAR/OUTBUF_GTS_AND ;
    wire \PAR/OFF/ASYNC_FF_GSR_OR ;
    wire \PAR/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[18]/SRNOT ;
    wire \AD[18]/IDELAY ;
    wire \AD[18]/OD ;
    wire \AD[18]/ENABLE ;
    wire \AD[18]/KEEPER ;
    wire \AD[18]/OUTBUF_GTS_AND ;
    wire \AD[18]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[18]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[18]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[12]/SRNOT ;
    wire \AD[12]/IDELAY ;
    wire \AD[12]/OD ;
    wire \AD[12]/ENABLE ;
    wire \AD[12]/KEEPER ;
    wire \AD[12]/OUTBUF_GTS_AND ;
    wire \AD[12]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[12]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[12]/TFF/ASYNC_FF_GSR_OR ;
    wire \CBE[1]/SRNOT ;
    wire \CBE[1]/IBUF ;
    wire \CBE[1]/IDELAY ;
    wire \CBE[1]/OD ;
    wire \CBE[1]/TNOT ;
    wire \CBE[1]/ENABLE ;
    wire \CBE[1]/KEEPER ;
    wire \CBE[1]/OUTBUF_GTS_AND ;
    wire \CBE[1]/IFF/ASYNC_FF_GSR_OR ;
    wire \CBE[1]/OFF/ASYNC_FF_GSR_OR ;
    wire \CBE[1]/TFF/ASYNC_FF_GSR_OR ;
    wire \TRDY/SRNOT ;
    wire \TRDY/IBUF ;
    wire \TRDY/IDELAY ;
    wire TRDY_out;
    wire \TRDY/TNOT ;
    wire TRDY_en;
    wire \TRDY/ENABLE ;
    wire \TRDY/KEEPER ;
    wire \TRDY/OUTBUF_GTS_AND ;
    wire \TRDY/IFF/ASYNC_FF_GSR_OR ;
    wire \TRDY/OFF/ASYNC_FF_GSR_OR ;
    wire \TRDY/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[11]/SRNOT ;
    wire \AD[11]/IDELAY ;
    wire \AD[11]/OD ;
    wire \AD[11]/ENABLE ;
    wire \AD[11]/KEEPER ;
    wire \AD[11]/OUTBUF_GTS_AND ;
    wire \AD[11]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[11]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[11]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[15]/SRNOT ;
    wire \AD[15]/IDELAY ;
    wire \AD[15]/OD ;
    wire \AD[15]/ENABLE ;
    wire \AD[15]/KEEPER ;
    wire \AD[15]/OUTBUF_GTS_AND ;
    wire \AD[15]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[15]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[15]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[14]/SRNOT ;
    wire \AD[14]/IDELAY ;
    wire \AD[14]/OD ;
    wire \AD[14]/ENABLE ;
    wire \AD[14]/KEEPER ;
    wire \AD[14]/OUTBUF_GTS_AND ;
    wire \AD[14]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[14]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[14]/TFF/ASYNC_FF_GSR_OR ;
    wire \DEVSEL/SRNOT ;
    wire \DEVSEL/IBUF ;
    wire \DEVSEL/IDELAY ;
    wire DEVSEL_out;
    wire \DEVSEL/TNOT ;
    wire DEVSEL_en;
    wire \DEVSEL/ENABLE ;
    wire \DEVSEL/KEEPER ;
    wire \DEVSEL/OUTBUF_GTS_AND ;
    wire \DEVSEL/IFF/ASYNC_FF_GSR_OR ;
    wire \DEVSEL/OFF/ASYNC_FF_GSR_OR ;
    wire \DEVSEL/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[10]/SRNOT ;
    wire \AD[10]/IDELAY ;
    wire \AD[10]/OD ;
    wire \AD[10]/ENABLE ;
    wire \AD[10]/KEEPER ;
    wire \AD[10]/OUTBUF_GTS_AND ;
    wire \AD[10]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[10]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[10]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[3]/SRNOT ;
    wire \AD[3]/IDELAY ;
    wire \AD[3]/OD ;
    wire \AD[3]/ENABLE ;
    wire \AD[3]/KEEPER ;
    wire \AD[3]/OUTBUF_GTS_AND ;
    wire \AD[3]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[3]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[3]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[9]/SRNOT ;
    wire \AD[9]/IDELAY ;
    wire \AD[9]/OD ;
    wire \AD[9]/ENABLE ;
    wire \AD[9]/KEEPER ;
    wire \AD[9]/OUTBUF_GTS_AND ;
    wire \AD[9]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[9]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[9]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[2]/SRNOT ;
    wire \AD[2]/IDELAY ;
    wire \AD[2]/OD ;
    wire \AD[2]/ENABLE ;
    wire \AD[2]/KEEPER ;
    wire \AD[2]/OUTBUF_GTS_AND ;
    wire \AD[2]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[2]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[2]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[8]/SRNOT ;
    wire \AD[8]/IDELAY ;
    wire \AD[8]/OD ;
    wire \AD[8]/ENABLE ;
    wire \AD[8]/KEEPER ;
    wire \AD[8]/OUTBUF_GTS_AND ;
    wire \AD[8]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[8]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[8]/TFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[29]/SRNOT ;
    wire \bridge/pci_target_unit/del_sync_addr_out[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync_addr_out[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \AD[1]/SRNOT ;
    wire \AD[1]/IDELAY ;
    wire \AD[1]/ENABLE ;
    wire \AD[1]/KEEPER ;
    wire \AD[1]/OUTBUF_GTS_AND ;
    wire \AD[1]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[1]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[1]/TFF/ASYNC_FF_GSR_OR ;
    wire \CBE[0]/SRNOT ;
    wire \CBE[0]/IBUF ;
    wire \CBE[0]/IDELAY ;
    wire \CBE[0]/OD ;
    wire \CBE[0]/TNOT ;
    wire \CBE[0]/ENABLE ;
    wire \CBE[0]/KEEPER ;
    wire \CBE[0]/OUTBUF_GTS_AND ;
    wire \CBE[0]/IFF/ASYNC_FF_GSR_OR ;
    wire \CBE[0]/OFF/ASYNC_FF_GSR_OR ;
    wire \CBE[0]/TFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[31]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \AD[6]/SRNOT ;
    wire \AD[6]/IDELAY ;
    wire \AD[6]/OD ;
    wire \AD[6]/ENABLE ;
    wire \AD[6]/KEEPER ;
    wire \AD[6]/OUTBUF_GTS_AND ;
    wire \AD[6]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[6]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[6]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[7]/SRNOT ;
    wire \AD[7]/IDELAY ;
    wire \AD[7]/OD ;
    wire \AD[7]/ENABLE ;
    wire \AD[7]/KEEPER ;
    wire \AD[7]/OUTBUF_GTS_AND ;
    wire \AD[7]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[7]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[7]/TFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[23]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \AD[5]/SRNOT ;
    wire \AD[5]/IDELAY ;
    wire \AD[5]/OD ;
    wire \AD[5]/ENABLE ;
    wire \AD[5]/KEEPER ;
    wire \AD[5]/OUTBUF_GTS_AND ;
    wire \AD[5]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[5]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[5]/TFF/ASYNC_FF_GSR_OR ;
    wire \GNT/IBUF ;
    wire \GNT/KEEPER ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[15]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \HSYNC/SRNOT ;
    wire \HSYNC/OD ;
    wire N_HSYNC;
    wire \HSYNC/KEEPER ;
    wire \HSYNC/OUTBUF_GTS_TRI ;
    wire \HSYNC/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[4]/SRNOT ;
    wire \AD[4]/IDELAY ;
    wire \AD[4]/OD ;
    wire \AD[4]/ENABLE ;
    wire \AD[4]/KEEPER ;
    wire \AD[4]/OUTBUF_GTS_AND ;
    wire \AD[4]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[4]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[4]/TFF/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[31]/SRNOT ;
    wire \CRT/pix_start_addr[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \REQ/SRNOT ;
    wire \REQ/OD ;
    wire REQ_out;
    wire \REQ/LOGIC_ZERO ;
    wire REQ_en;
    wire \REQ/ENABLE ;
    wire \REQ/KEEPER ;
    wire \REQ/OUTBUF_GTS_AND ;
    wire \REQ/OFF/ASYNC_FF_GSR_OR ;
    wire \REQ/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[0]/SRNOT ;
    wire \AD[0]/IDELAY ;
    wire \AD[0]/OD ;
    wire \AD[0]/ENABLE ;
    wire \AD[0]/KEEPER ;
    wire \AD[0]/OUTBUF_GTS_AND ;
    wire \AD[0]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[0]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[0]/TFF/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[23]/SRNOT ;
    wire \CRT/pix_start_addr[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \VSYNC/SRNOT ;
    wire \VSYNC/OD ;
    wire N_VSYNC;
    wire \VSYNC/KEEPER ;
    wire \VSYNC/OUTBUF_GTS_TRI ;
    wire \VSYNC/OFF/ASYNC_FF_GSR_OR ;
    wire \LED/OD ;
    wire \LED/KEEPER ;
    wire \LED/OUTBUF_GTS_TRI ;
    wire \CRT/pix_start_addr[15]/SRNOT ;
    wire \CRT/pix_start_addr[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \AD[31]/SRNOT ;
    wire \AD[31]/IDELAY ;
    wire \AD[31]/ENABLE ;
    wire \AD[31]/KEEPER ;
    wire \AD[31]/OUTBUF_GTS_AND ;
    wire \AD[31]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[31]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[31]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[30]/SRNOT ;
    wire \AD[30]/IDELAY ;
    wire \AD[30]/ENABLE ;
    wire \AD[30]/KEEPER ;
    wire \AD[30]/OUTBUF_GTS_AND ;
    wire \AD[30]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[30]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[30]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[29]/SRNOT ;
    wire \AD[29]/IDELAY ;
    wire \AD[29]/OD ;
    wire \AD[29]/ENABLE ;
    wire \AD[29]/KEEPER ;
    wire \AD[29]/OUTBUF_GTS_AND ;
    wire \AD[29]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[29]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[29]/TFF/ASYNC_FF_GSR_OR ;
    wire \AD[28]/SRNOT ;
    wire \AD[28]/IDELAY ;
    wire \AD[28]/OD ;
    wire \AD[28]/ENABLE ;
    wire \AD[28]/KEEPER ;
    wire \AD[28]/OUTBUF_GTS_AND ;
    wire \AD[28]/IFF/ASYNC_FF_GSR_OR ;
    wire \AD[28]/OFF/ASYNC_FF_GSR_OR ;
    wire \AD[28]/TFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_bc_out[1]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_bc_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_bc_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \RGB[14]/SRNOT ;
    wire \RGB[14]/OD ;
    wire \RGB[14]/KEEPER ;
    wire \RGB[14]/OUTBUF_GTS_TRI ;
    wire \RGB[14]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[7]/SRNOT ;
    wire \RGB[7]/KEEPER ;
    wire \RGB[7]/OUTBUF_GTS_TRI ;
    wire \RGB[7]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[15]/SRNOT ;
    wire \RGB[15]/OD ;
    wire \RGB[15]/KEEPER ;
    wire \RGB[15]/OUTBUF_GTS_TRI ;
    wire \RGB[15]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[8]/SRNOT ;
    wire \RGB[8]/OD ;
    wire \RGB[8]/KEEPER ;
    wire \RGB[8]/OUTBUF_GTS_TRI ;
    wire \RGB[8]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[9]/SRNOT ;
    wire \RGB[9]/OD ;
    wire \RGB[9]/KEEPER ;
    wire \RGB[9]/OUTBUF_GTS_TRI ;
    wire \RGB[9]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[4]/SRNOT ;
    wire \RGB[4]/OD ;
    wire \RGB[4]/KEEPER ;
    wire \RGB[4]/OUTBUF_GTS_TRI ;
    wire \RGB[4]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[5]/SRNOT ;
    wire \RGB[5]/OD ;
    wire \RGB[5]/KEEPER ;
    wire \RGB[5]/OUTBUF_GTS_TRI ;
    wire \RGB[5]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[10]/SRNOT ;
    wire \RGB[10]/OD ;
    wire \RGB[10]/KEEPER ;
    wire \RGB[10]/OUTBUF_GTS_TRI ;
    wire \RGB[10]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[6]/SRNOT ;
    wire \RGB[6]/KEEPER ;
    wire \RGB[6]/OUTBUF_GTS_TRI ;
    wire \RGB[6]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[11]/SRNOT ;
    wire \RGB[11]/OD ;
    wire \RGB[11]/KEEPER ;
    wire \RGB[11]/OUTBUF_GTS_TRI ;
    wire \RGB[11]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[12]/SRNOT ;
    wire \RGB[12]/OD ;
    wire \RGB[12]/KEEPER ;
    wire \RGB[12]/OUTBUF_GTS_TRI ;
    wire \RGB[12]/OFF/ASYNC_FF_GSR_OR ;
    wire \RGB[13]/SRNOT ;
    wire \RGB[13]/OD ;
    wire \RGB[13]/KEEPER ;
    wire \RGB[13]/OUTBUF_GTS_TRI ;
    wire \RGB[13]/OFF/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[25]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[17]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[25]/SRNOT ;
    wire \CRT/pix_start_addr[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[17]/SRNOT ;
    wire \CRT/pix_start_addr[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_bc_out[3]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_bc_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_bc_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pci_target_if/C5316/C2/N8 ;
    wire \bridge/pci_target_unit/pci_target_if/N5157/F5MUX ;
    wire \bridge/pci_target_unit/pci_target_if/C5316/C2/N7 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ONE ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3384/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C3/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3384/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3384/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3384/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3384/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3386/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C5/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3386/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3386/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3386/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3386/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3386/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3388/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C7/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3388/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3388/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3388/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3388/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3388/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3390/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C9/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3390/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3390/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3390/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3390/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3390/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3392/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C11/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3392/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3392/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3392/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3392/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3392/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3394/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C13/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3394/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3394/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3394/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3394/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3394/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[27]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3396/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C15/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3396/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3396/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3396/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3396/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3396/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[19]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3398/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C17/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3398/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3398/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3398/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3398/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3398/XORF ;
    wire \CRT/pix_start_addr[27]/SRNOT ;
    wire \CRT/pix_start_addr[27]/FROM ;
    wire \CRT/pix_start_addr[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3400/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C19/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3400/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3400/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3400/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3400/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3400/XORF ;
    wire \CRT/pix_start_addr[19]/SRNOT ;
    wire \CRT/pix_start_addr[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3402/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C21/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3402/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3402/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3402/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3402/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3402/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3404/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C23/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3404/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3404/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3404/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3404/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3404/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3406/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C25/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3406/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3406/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3406/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3406/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3406/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3408/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C27/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3408/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3408/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3408/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3408/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3408/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3410/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C29/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3410/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3410/CYMUXG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3410/GROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3410/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3410/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[29]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3412/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C31/C1/O ;
    wire \bridge/wishbone_slave_unit/pcim_if_address_out[31]_rt ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3412/FROM ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3412/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3412/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/N738/LOGIC_ONE ;
    wire \CRT/ssvga_fifo/N738/XORG ;
    wire \CRT/ssvga_fifo/C748/C3/C1/O ;
    wire \CRT/ssvga_fifo/N738/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/N738/CYMUXG ;
    wire \CRT/ssvga_fifo/N738/GROM ;
    wire \CRT/ssvga_fifo/N738/FROM ;
    wire \CRT/ssvga_fifo/N738/XORF ;
    wire \CRT/pix_start_addr[29]/SRNOT ;
    wire \CRT/pix_start_addr[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/pix_start_addr[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/N740/XORG ;
    wire \CRT/ssvga_fifo/C748/C5/C1/O ;
    wire \CRT/ssvga_fifo/N740/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/N740/CYMUXG ;
    wire \CRT/ssvga_fifo/N740/GROM ;
    wire \CRT/ssvga_fifo/N740/FROM ;
    wire \CRT/ssvga_fifo/N740/XORF ;
    wire \CRT/ssvga_fifo/N742/XORG ;
    wire \CRT/ssvga_fifo/C748/C7/C1/O ;
    wire \CRT/ssvga_fifo/N742/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/N742/CYMUXG ;
    wire \CRT/ssvga_fifo/N742/GROM ;
    wire \CRT/ssvga_fifo/N742/FROM ;
    wire \CRT/ssvga_fifo/N742/XORF ;
    wire \CRT/ssvga_fifo/N744/XORG ;
    wire \CRT/ssvga_fifo/C748/C9/C1/O ;
    wire \CRT/ssvga_fifo/N744/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/N744/CYMUXG ;
    wire \CRT/ssvga_fifo/N744/GROM ;
    wire \CRT/ssvga_fifo/N744/FROM ;
    wire \CRT/ssvga_fifo/N744/XORF ;
    wire \bridge/configuration/pci_error_rty_exp_set/LOGIC_ONE ;
    wire \bridge/configuration/pci_error_rty_exp_set/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/N746/XORG ;
    wire \CRT/ssvga_fifo/C748/C11/C1/O ;
    wire \CRT/ssvga_fifo/rd_ptr_plus1[9]_rt ;
    wire \CRT/ssvga_fifo/N746/FROM ;
    wire \CRT/ssvga_fifo/N746/XORF ;
    wire \CRT/ssvga_fifo/N746/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1515/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1515/XORG ;
    wire \CRT/ssvga_wbm_if/C1472/C3/C1/O ;
    wire \CRT/ssvga_wbm_if/N1515/CYMUXG ;
    wire N12625;
    wire N12642;
    wire \CRT/ssvga_wbm_if/N1515/XORF ;
    wire \bridge/pci_target_unit/pci_target_if/bckp_trdy_reg/SRNOT ;
    wire \bridge/pci_target_unit/pci_target_if/bckp_trdy_reg/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1517/XORG ;
    wire \CRT/ssvga_wbm_if/C1472/C5/C1/O ;
    wire \CRT/ssvga_wbm_if/N1517/CYMUXG ;
    wire N12619;
    wire N12650;
    wire \CRT/ssvga_wbm_if/N1517/XORF ;
    wire \bridge/conf_cache_line_size_out[1]/SRNOT ;
    wire \bridge/conf_cache_line_size_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_cache_line_size_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1519/XORG ;
    wire \CRT/ssvga_wbm_if/C1472/C7/C1/O ;
    wire \CRT/ssvga_wbm_if/N1519/CYMUXG ;
    wire N12623;
    wire N12646;
    wire \CRT/ssvga_wbm_if/N1519/XORF ;
    wire \CRT/ssvga_wbm_if/N1521/XORG ;
    wire \CRT/ssvga_wbm_if/C1472/C9/C1/O ;
    wire \CRT/ssvga_wbm_if/N1521/CYMUXG ;
    wire N12621;
    wire N12648;
    wire \CRT/ssvga_wbm_if/N1521/XORF ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1523/XORG ;
    wire \CRT/ssvga_wbm_if/C1472/C11/C1/O ;
    wire \CRT/ssvga_wbm_if/N1523/CYMUXG ;
    wire N12644;
    wire N12627;
    wire \CRT/ssvga_wbm_if/N1523/XORF ;
    wire \bridge/conf_cache_line_size_out[3]/SRNOT ;
    wire \bridge/conf_cache_line_size_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_cache_line_size_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1525/XORG ;
    wire \CRT/ssvga_wbm_if/C1472/C13/C1/O ;
    wire \CRT/ssvga_wbm_if/N1525/CYMUXG ;
    wire N12631;
    wire N12638;
    wire \CRT/ssvga_wbm_if/N1525/XORF ;
    wire \CRT/ssvga_wbm_if/N1527/XORG ;
    wire \CRT/ssvga_wbm_if/C1472/C15/C1/O ;
    wire \CRT/ssvga_wbm_if/N1527/CYMUXG ;
    wire N12633;
    wire N12636;
    wire \CRT/ssvga_wbm_if/N1527/XORF ;
    wire \CRT/ssvga_wbm_if/N1529/XORG ;
    wire \CRT/ssvga_wbm_if/C1472/C17/C1/O ;
    wire \CRT/ssvga_wbm_if/N1529/CYMUXG ;
    wire N12629;
    wire N12640;
    wire \CRT/ssvga_wbm_if/N1529/XORF ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/N800/LOGIC_ONE ;
    wire \CRT/ssvga_fifo/N800/XORG ;
    wire \CRT/ssvga_fifo/C749/C3/C1/O ;
    wire \CRT/ssvga_fifo/N800/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/N800/CYMUXG ;
    wire \CRT/ssvga_fifo/N800/GROM ;
    wire \CRT/ssvga_fifo/N800/FROM ;
    wire \CRT/ssvga_fifo/N800/XORF ;
    wire \bridge/conf_cache_line_size_out[5]/SRNOT ;
    wire \bridge/conf_cache_line_size_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_cache_line_size_out[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_fifo/N802/XORG ;
    wire \CRT/ssvga_fifo/C749/C5/C1/O ;
    wire \CRT/ssvga_fifo/N802/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/N802/CYMUXG ;
    wire \CRT/ssvga_fifo/N802/GROM ;
    wire \CRT/ssvga_fifo/N802/FROM ;
    wire \CRT/ssvga_fifo/N802/XORF ;
    wire \CRT/ssvga_fifo/N804/XORG ;
    wire \CRT/ssvga_fifo/C749/C7/C1/O ;
    wire \CRT/ssvga_fifo/N804/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/N804/CYMUXG ;
    wire \CRT/ssvga_fifo/N804/GROM ;
    wire \CRT/ssvga_fifo/N804/FROM ;
    wire \CRT/ssvga_fifo/N804/XORF ;
    wire \CRT/ssvga_fifo/N806/XORG ;
    wire \CRT/ssvga_fifo/C749/C9/C1/O ;
    wire \CRT/ssvga_fifo/wr_ptr_plus1[7]_rt ;
    wire \CRT/ssvga_fifo/N806/FROM ;
    wire \CRT/ssvga_fifo/N806/XORF ;
    wire \CRT/ssvga_fifo/N806/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[4]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/N1235/LOGIC_ONE ;
    wire \bridge/pci_target_unit/del_sync/N1235/XORG ;
    wire \bridge/pci_target_unit/del_sync/C1264/C3/C1/O ;
    wire \bridge/pci_target_unit/del_sync/N1235/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/del_sync/N1235/CYMUXG ;
    wire \bridge/pci_target_unit/del_sync/N1235/GROM ;
    wire \bridge/pci_target_unit/del_sync/N1235/FROM ;
    wire \bridge/pci_target_unit/del_sync/N1235/XORF ;
    wire \bridge/conf_cache_line_size_out[7]/SRNOT ;
    wire \bridge/conf_cache_line_size_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/conf_cache_line_size_out[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/N1237/XORG ;
    wire \bridge/pci_target_unit/del_sync/C1264/C5/C1/O ;
    wire \bridge/pci_target_unit/del_sync/N1237/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/del_sync/N1237/CYMUXG ;
    wire \bridge/pci_target_unit/del_sync/N1237/GROM ;
    wire \bridge/pci_target_unit/del_sync/N1237/FROM ;
    wire \bridge/pci_target_unit/del_sync/N1237/XORF ;
    wire \bridge/pci_target_unit/del_sync/N1239/XORG ;
    wire \bridge/pci_target_unit/del_sync/C1264/C7/C1/O ;
    wire \bridge/pci_target_unit/del_sync/N1239/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/del_sync/N1239/CYMUXG ;
    wire \bridge/pci_target_unit/del_sync/N1239/GROM ;
    wire \bridge/pci_target_unit/del_sync/N1239/FROM ;
    wire \bridge/pci_target_unit/del_sync/N1239/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[1]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/N1241/XORG ;
    wire \bridge/pci_target_unit/del_sync/C1264/C9/C1/O ;
    wire \bridge/pci_target_unit/del_sync/N1241/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/del_sync/N1241/CYMUXG ;
    wire \bridge/pci_target_unit/del_sync/N1241/GROM ;
    wire \bridge/pci_target_unit/del_sync/N1241/FROM ;
    wire \bridge/pci_target_unit/del_sync/N1241/XORF ;
    wire \bridge/pci_target_unit/del_sync/N1243/XORG ;
    wire \bridge/pci_target_unit/del_sync/C1264/C11/C1/O ;
    wire \bridge/pci_target_unit/del_sync/N1243/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/del_sync/N1243/CYMUXG ;
    wire \bridge/pci_target_unit/del_sync/N1243/GROM ;
    wire \bridge/pci_target_unit/del_sync/N1243/FROM ;
    wire \bridge/pci_target_unit/del_sync/N1243/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[3]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/N1245/XORG ;
    wire \bridge/pci_target_unit/del_sync/C1264/C13/C1/O ;
    wire \bridge/pci_target_unit/del_sync/N1245/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/del_sync/N1245/CYMUXG ;
    wire \bridge/pci_target_unit/del_sync/N1245/GROM ;
    wire \bridge/pci_target_unit/del_sync/N1245/FROM ;
    wire \bridge/pci_target_unit/del_sync/N1245/XORF ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/BYNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/SRNOT ;
    wire \bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/N1247/XORG ;
    wire \bridge/pci_target_unit/del_sync/C1264/C15/C1/O ;
    wire \bridge/pci_target_unit/del_sync/N1247/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/del_sync/N1247/CYMUXG ;
    wire \bridge/pci_target_unit/del_sync/N1247/GROM ;
    wire \bridge/pci_target_unit/del_sync/N1247/FROM ;
    wire \bridge/pci_target_unit/del_sync/N1247/XORF ;
    wire \bridge/pci_target_unit/del_sync/N1249/XORG ;
    wire \bridge/pci_target_unit/del_sync/C1264/C17/C1/O ;
    wire \bridge/pci_target_unit/del_sync/N1249/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/del_sync/N1249/CYMUXG ;
    wire \bridge/pci_target_unit/del_sync/N1249/GROM ;
    wire \bridge/pci_target_unit/del_sync/N1249/FROM ;
    wire \bridge/pci_target_unit/del_sync/N1249/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[5]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/del_sync/comp_cycle_count[16]_rt ;
    wire \bridge/pci_target_unit/del_sync/N1251/XORF ;
    wire \CRT/ssvga_wbm_if/N1717/LOGIC_ONE ;
    wire \CRT/ssvga_wbm_if/N1717/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C3/C1/O ;
    wire \CRT/ssvga_wbm_if/N1717/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1717/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1717/GROM ;
    wire \CRT/ssvga_wbm_if/N1717/FROM ;
    wire \CRT/ssvga_wbm_if/N1717/XORF ;
    wire \CRT/ssvga_wbm_if/N1719/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C5/C1/O ;
    wire \CRT/ssvga_wbm_if/N1719/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1719/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1719/GROM ;
    wire \CRT/ssvga_wbm_if/N1719/FROM ;
    wire \CRT/ssvga_wbm_if/N1719/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[7]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1721/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C7/C1/O ;
    wire \CRT/ssvga_wbm_if/N1721/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1721/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1721/GROM ;
    wire \CRT/ssvga_wbm_if/N1721/FROM ;
    wire \CRT/ssvga_wbm_if/N1721/XORF ;
    wire \CRT/ssvga_wbm_if/N1723/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C9/C1/O ;
    wire \CRT/ssvga_wbm_if/N1723/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1723/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1723/GROM ;
    wire \CRT/ssvga_wbm_if/N1723/FROM ;
    wire \CRT/ssvga_wbm_if/N1723/XORF ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[9]/SRNOT ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[9]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/pcit_if_addr_out[9]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1725/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C11/C1/O ;
    wire \CRT/ssvga_wbm_if/N1725/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1725/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1725/GROM ;
    wire \CRT/ssvga_wbm_if/N1725/FROM ;
    wire \CRT/ssvga_wbm_if/N1725/XORF ;
    wire \CRT/ssvga_wbm_if/N1727/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C13/C1/O ;
    wire \CRT/ssvga_wbm_if/N1727/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1727/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1727/GROM ;
    wire \CRT/ssvga_wbm_if/N1727/FROM ;
    wire \CRT/ssvga_wbm_if/N1727/XORF ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[4]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1729/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C15/C1/O ;
    wire \CRT/ssvga_wbm_if/N1729/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1729/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1729/GROM ;
    wire \CRT/ssvga_wbm_if/N1729/FROM ;
    wire \CRT/ssvga_wbm_if/N1729/XORF ;
    wire \bridge/out_bckp_irdy_en_out/SRNOT ;
    wire \bridge/out_bckp_irdy_en_out/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1731/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C17/C1/O ;
    wire \CRT/ssvga_wbm_if/N1731/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1731/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1731/GROM ;
    wire \CRT/ssvga_wbm_if/N1731/FROM ;
    wire \CRT/ssvga_wbm_if/N1731/XORF ;
    wire \CRT/ssvga_wbm_if/N1733/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C19/C1/O ;
    wire \CRT/ssvga_wbm_if/N1733/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1733/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1733/GROM ;
    wire \CRT/ssvga_wbm_if/N1733/FROM ;
    wire \CRT/ssvga_wbm_if/N1733/XORF ;
    wire \bridge/parity_checker/check_perr/SRNOT ;
    wire \bridge/parity_checker/check_perr/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1735/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C21/C1/O ;
    wire \CRT/ssvga_wbm_if/N1735/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1735/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1735/GROM ;
    wire \CRT/ssvga_wbm_if/N1735/FROM ;
    wire \CRT/ssvga_wbm_if/N1735/XORF ;
    wire \bridge/pci_target_unit/del_sync/sync_comp_req_pending/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/sync_comp_req_pending/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1737/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C23/C1/O ;
    wire \CRT/ssvga_wbm_if/N1737/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1737/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1737/GROM ;
    wire \CRT/ssvga_wbm_if/N1737/FROM ;
    wire \CRT/ssvga_wbm_if/N1737/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1739/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C25/C1/O ;
    wire \CRT/ssvga_wbm_if/N1739/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1739/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1739/GROM ;
    wire \CRT/ssvga_wbm_if/N1739/FROM ;
    wire \CRT/ssvga_wbm_if/N1739/XORF ;
    wire \crt_vsync/BYNOT ;
    wire \crt_vsync/SRNOT ;
    wire \crt_vsync/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1741/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C27/C1/O ;
    wire \CRT/ssvga_wbm_if/N1741/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1741/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1741/GROM ;
    wire \CRT/ssvga_wbm_if/N1741/FROM ;
    wire \CRT/ssvga_wbm_if/N1741/XORF ;
    wire \bridge/conf_perr_response_out/SRNOT ;
    wire \bridge/conf_perr_response_out/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1743/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C29/C1/O ;
    wire \CRT/ssvga_wbm_if/N1743/LOGIC_ZERO ;
    wire \CRT/ssvga_wbm_if/N1743/CYMUXG ;
    wire \CRT/ssvga_wbm_if/N1743/GROM ;
    wire \CRT/ssvga_wbm_if/N1743/FROM ;
    wire \CRT/ssvga_wbm_if/N1743/XORF ;
    wire \bridge/pci_target_unit/del_sync/comp_done_reg_main/SRNOT ;
    wire \bridge/pci_target_unit/del_sync/comp_done_reg_main/FFY/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_wbm_if/N1745/XORG ;
    wire \CRT/ssvga_wbm_if/C1473/C31/C1/O ;
    wire \bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]_rt ;
    wire \CRT/ssvga_wbm_if/N1745/FROM ;
    wire \CRT/ssvga_wbm_if/N1745/XORF ;
    wire \CRT/ssvga_wbm_if/N1745/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N326/LOGIC_ONE ;
    wire \CRT/ssvga_crtc/N326/XORG ;
    wire \CRT/ssvga_crtc/C529/C3/C1/O ;
    wire \CRT/ssvga_crtc/N326/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N326/CYMUXG ;
    wire \CRT/ssvga_crtc/N326/GROM ;
    wire \CRT/ssvga_crtc/N326/FROM ;
    wire \CRT/ssvga_crtc/N326/XORF ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/N328/XORG ;
    wire \CRT/ssvga_crtc/C529/C5/C1/O ;
    wire \CRT/ssvga_crtc/N328/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N328/CYMUXG ;
    wire \CRT/ssvga_crtc/N328/GROM ;
    wire \CRT/ssvga_crtc/N328/FROM ;
    wire \CRT/ssvga_crtc/N328/XORF ;
    wire \CRT/ssvga_crtc/N330/XORG ;
    wire \CRT/ssvga_crtc/C529/C7/C1/O ;
    wire \CRT/ssvga_crtc/N330/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N330/CYMUXG ;
    wire \CRT/ssvga_crtc/N330/GROM ;
    wire \CRT/ssvga_crtc/N330/FROM ;
    wire \CRT/ssvga_crtc/N330/XORF ;
    wire \N12322/GROM ;
    wire \N12322/FROM ;
    wire \CRT/ssvga_crtc/N332/XORG ;
    wire \CRT/ssvga_crtc/C529/C9/C1/O ;
    wire \CRT/ssvga_crtc/N332/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N332/CYMUXG ;
    wire \CRT/ssvga_crtc/N332/GROM ;
    wire \CRT/ssvga_crtc/N332/FROM ;
    wire \CRT/ssvga_crtc/N332/XORF ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFY/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFX/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \CRT/ssvga_crtc/N334/XORG ;
    wire \CRT/ssvga_crtc/C529/C11/C1/O ;
    wire \CRT/ssvga_crtc/vcntr[9]_rt ;
    wire \CRT/ssvga_crtc/N334/FROM ;
    wire \CRT/ssvga_crtc/N334/XORF ;
    wire \CRT/ssvga_crtc/N334/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ONE ;
    wire \bridge/pci_target_unit/wishbone_master/N3068/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3410/C3/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/wishbone_master/N3068/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/C3413/N12 ;
    wire \bridge/pci_target_unit/wishbone_master/C3413/N6 ;
    wire \bridge/pci_target_unit/wishbone_master/N3068/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3070/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3410/C5/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3070/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/wishbone_master/N3070/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/C3413/N24 ;
    wire \bridge/pci_target_unit/wishbone_master/C3413/N18 ;
    wire \bridge/pci_target_unit/wishbone_master/N3070/XORF ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[4]/FFY/SET ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/N3072/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3410/C7/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3072/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/wishbone_master/N3072/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/C3413/N36 ;
    wire \bridge/pci_target_unit/wishbone_master/C3413/N30 ;
    wire \bridge/pci_target_unit/wishbone_master/N3072/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3074/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3410/C9/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/C3413/N48 ;
    wire \bridge/pci_target_unit/wishbone_master/C3413/N42 ;
    wire \bridge/pci_target_unit/wishbone_master/N3074/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3074/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync_comp_flush_out/SRNOT ;
    wire \bridge/wishbone_slave_unit/del_sync_comp_flush_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/N2983/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/wishbone_master/N2983/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C2/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2983/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2983/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2983/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2983/XORF ;
    wire \bridge/conf_serr_enable_out/SRNOT ;
    wire \bridge/conf_serr_enable_out/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/N2985/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C4/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2985/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2985/GROM ;
    wire N12692;
    wire \bridge/pci_target_unit/wishbone_master/N2985/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N2987/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C6/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2987/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2987/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2987/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2987/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N2989/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C8/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2989/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2989/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2989/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2989/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N2991/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C10/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2991/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2991/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2991/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2991/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N2993/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C12/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2993/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2993/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2993/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2993/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N2995/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C14/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2995/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2995/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2995/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2995/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N2997/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C16/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2997/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2997/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2997/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2997/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N2999/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C18/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N2999/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N2999/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2999/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N2999/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3001/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C20/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3001/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N3001/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3001/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3001/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3003/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C22/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3003/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N3003/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3003/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3003/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3005/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C24/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3005/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N3005/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3005/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3005/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3007/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C26/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3007/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N3007/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3007/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3007/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3009/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C28/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3009/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N3009/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3009/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3009/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3011/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C30/C2/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3011/CYMUXG ;
    wire \bridge/pci_target_unit/wishbone_master/N3011/GROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3011/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3011/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3013/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3409/C32/C2/O ;
    wire \bridge/pciu_err_addr_out[31]_rt ;
    wire \bridge/pci_target_unit/wishbone_master/N3013/FROM ;
    wire \bridge/pci_target_unit/wishbone_master/N3013/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3110/LOGIC_ZERO ;
    wire \bridge/pci_target_unit/wishbone_master/N3110/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3411/C3/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3110/CYMUXG ;
    wire N12696;
    wire N12694;
    wire \bridge/pci_target_unit/wishbone_master/N3110/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3112/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3411/C5/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3112/CYMUXG ;
    wire N12700;
    wire N12698;
    wire \bridge/pci_target_unit/wishbone_master/N3112/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3114/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3411/C7/C1/O ;
    wire \bridge/pci_target_unit/wishbone_master/N3114/CYMUXG ;
    wire N12704;
    wire N12702;
    wire \bridge/pci_target_unit/wishbone_master/N3114/XORF ;
    wire \bridge/pci_target_unit/wishbone_master/N3116/XORG ;
    wire \bridge/pci_target_unit/wishbone_master/C3411/C9/C1/O ;
    wire N12708;
    wire N12706;
    wire \bridge/pci_target_unit/wishbone_master/N3116/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2618/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2618/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C3/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2618/CYMUXG ;
    wire N12657;
    wire N12655;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2618/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2620/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C5/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2620/CYMUXG ;
    wire N12661;
    wire N12659;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2620/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2622/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C7/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2622/CYMUXG ;
    wire N12665;
    wire N12663;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2622/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2624/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C9/C1/O ;
    wire N12669;
    wire N12667;
    wire \bridge/wishbone_slave_unit/pci_initiator_sm/N2624/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ONE ;
    wire \bridge/wishbone_slave_unit/del_sync/N140/XORG ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C3/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync/N140/CYMUXG ;
    wire \bridge/wishbone_slave_unit/del_sync/N140/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N140/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N140/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/N142/XORG ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C5/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/N142/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync/N142/CYMUXG ;
    wire \bridge/wishbone_slave_unit/del_sync/N142/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N142/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N142/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/N144/XORG ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C7/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/N144/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync/N144/CYMUXG ;
    wire \bridge/wishbone_slave_unit/del_sync/N144/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N144/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N144/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/N146/XORG ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C9/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/N146/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync/N146/CYMUXG ;
    wire \bridge/wishbone_slave_unit/del_sync/N146/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N146/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N146/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/N148/XORG ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C11/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/N148/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync/N148/CYMUXG ;
    wire \bridge/wishbone_slave_unit/del_sync/N148/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N148/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N148/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/N150/XORG ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C13/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/N150/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync/N150/CYMUXG ;
    wire \bridge/wishbone_slave_unit/del_sync/N150/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N150/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N150/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/N152/XORG ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C15/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/N152/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync/N152/CYMUXG ;
    wire \bridge/wishbone_slave_unit/del_sync/N152/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N152/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N152/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/N154/XORG ;
    wire \bridge/wishbone_slave_unit/del_sync/C24/C17/C1/O ;
    wire \bridge/wishbone_slave_unit/del_sync/N154/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/del_sync/N154/CYMUXG ;
    wire \bridge/wishbone_slave_unit/del_sync/N154/GROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N154/FROM ;
    wire \bridge/wishbone_slave_unit/del_sync/N154/XORF ;
    wire \bridge/wishbone_slave_unit/del_sync/comp_cycle_count[16]_rt ;
    wire \bridge/wishbone_slave_unit/del_sync/N156/XORF ;
    wire \CRT/ssvga_crtc/N400/LOGIC_ONE ;
    wire \CRT/ssvga_crtc/N400/XORG ;
    wire \CRT/ssvga_crtc/C530/C3/C1/O ;
    wire \CRT/ssvga_crtc/N400/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N400/CYMUXG ;
    wire \CRT/ssvga_crtc/N400/GROM ;
    wire \CRT/ssvga_crtc/N400/FROM ;
    wire \CRT/ssvga_crtc/N400/XORF ;
    wire \CRT/ssvga_crtc/N402/XORG ;
    wire \CRT/ssvga_crtc/C530/C5/C1/O ;
    wire \CRT/ssvga_crtc/N402/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N402/CYMUXG ;
    wire \CRT/ssvga_crtc/N402/GROM ;
    wire \CRT/ssvga_crtc/N402/FROM ;
    wire \CRT/ssvga_crtc/N402/XORF ;
    wire \CRT/ssvga_crtc/N404/XORG ;
    wire \CRT/ssvga_crtc/C530/C7/C1/O ;
    wire \CRT/ssvga_crtc/N404/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N404/CYMUXG ;
    wire \CRT/ssvga_crtc/N404/GROM ;
    wire \CRT/ssvga_crtc/N404/FROM ;
    wire \CRT/ssvga_crtc/N404/XORF ;
    wire \CRT/ssvga_crtc/N406/XORG ;
    wire \CRT/ssvga_crtc/C530/C9/C1/O ;
    wire \CRT/ssvga_crtc/N406/LOGIC_ZERO ;
    wire \CRT/ssvga_crtc/N406/CYMUXG ;
    wire \CRT/ssvga_crtc/N406/GROM ;
    wire \CRT/ssvga_crtc/N406/FROM ;
    wire \CRT/ssvga_crtc/N406/XORF ;
    wire \CRT/ssvga_crtc/N408/XORG ;
    wire \CRT/ssvga_crtc/C530/C11/C1/O ;
    wire \CRT/ssvga_crtc/hcntr[9]_rt ;
    wire \CRT/ssvga_crtc/N408/FROM ;
    wire \CRT/ssvga_crtc/N408/XORF ;
    wire \CRT/ssvga_crtc/N408/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3190/LOGIC_ZERO ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3190/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C3/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3190/CYMUXG ;
    wire N12675;
    wire N12673;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3190/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3192/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C5/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3192/CYMUXG ;
    wire N12679;
    wire N12677;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3192/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3194/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C7/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3194/CYMUXG ;
    wire N12683;
    wire N12681;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3194/XORF ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3196/XORG ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C9/C1/O ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3196/CYMUXG ;
    wire N12687;
    wire N12685;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3196/XORF ;
    wire N12689;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/N3198/XORF ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[25]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[25]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[25]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[17]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[17]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[17]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N12 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N6 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N60 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N54 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N108 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N102 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[1]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3414/N6 ;
    wire \bridge/pci_target_unit/wishbone_master/C3414/N12 ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[27]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[27]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[27]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[19]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[19]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[19]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N48 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N42 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N96 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N90 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[3]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3414/N18 ;
    wire \bridge/pci_target_unit/wishbone_master/C3414/N24 ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[29]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[29]/GROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[29]/FROM ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pcim_if_data_out[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[1]/GROM ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[1]/FFY/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[1]/FFX/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_waddr[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N36 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N30 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N84 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N78 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[5]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3414/N30 ;
    wire \bridge/pci_target_unit/wishbone_master/C3414/N36 ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[5]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[5]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFY/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFX/RST ;
    wire \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/SRNOT ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N24 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/C13/N18 ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/mrl_en/SRNOT ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/mrl_en/GROM ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/mrl_en/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/wishbone_slave/mrl_en/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[7]/SRNOT ;
    wire \bridge/pci_target_unit/wishbone_master/C3414/N42 ;
    wire \bridge/pci_target_unit/wishbone_master/C3414/N48 ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[7]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/pci_target_unit/wishbone_master/cache_line[7]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/GROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty111 ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/FROM ;
    wire \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/outGreyCount[1]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/outGreyCount[1]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/outGreyCount[3]/SRNOT ;
    wire \bridge/wishbone_slave_unit/fifos/outGreyCount[3]/FFY/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/outGreyCount[3]/FFX/ASYNC_FF_GSR_OR ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_1/LOGIC_ONE ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_1/RSTANOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_1/RSTBNOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_1/WEANOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_1/INT_SIG ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_2/LOGIC_ONE ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_2/RSTANOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_2/RSTBNOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_2/WEANOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_2/INT_SIG ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA0 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA1 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA2 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA3 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA4 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA5 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA6 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA7 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA8 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA9 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA10 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA11 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA14 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA15 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB4 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB5 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB6 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB7 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB8 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB9 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB10 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB11 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB13 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB14 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB15 ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/LOGIC_ONE ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/RSTANOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/RSTBNOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/WEANOT ;
    wire \bridge/wishbone_slave_unit/fifos/dpram16_3/INT_SIG ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB0 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB1 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB2 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB3 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB4 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB5 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB6 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB7 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB8 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB9 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB10 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB11 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB12 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB13 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB14 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/DOB15 ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ONE ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/RSTANOT ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/RSTBNOT ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/ramb4_s8_0/INT_SIG ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB0 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB1 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB2 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB3 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB4 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB5 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB6 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB7 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB8 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB9 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB10 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB11 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB12 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB13 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB14 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/DOB15 ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ONE ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/RSTANOT ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/RSTBNOT ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ZERO ;
    wire \CRT/ssvga_fifo/ramb4_s8_1/INT_SIG ;
    wire \CRT/ssvga_pallete/DOB0 ;
    wire \CRT/ssvga_pallete/DOB1 ;
    wire \CRT/ssvga_pallete/DOB2 ;
    wire \CRT/ssvga_pallete/DOB3 ;
    wire \CRT/ssvga_pallete/LOGIC_ONE ;
    wire \CRT/ssvga_pallete/RSTANOT ;
    wire \CRT/ssvga_pallete/RSTBNOT ;
    wire \CRT/ssvga_pallete/LOGIC_ZERO ;
    wire \CRT/ssvga_pallete/INT_SIG ;
    wire \bridge/pci_target_unit/fifos/dpram16_1/RSTANOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_1/RSTBNOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_1/WEANOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_1/INT_SIG ;
    wire \bridge/pci_target_unit/fifos/dpram16_2/RSTANOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_2/RSTBNOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_2/WEANOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_2/INT_SIG ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA0 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA1 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA2 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA3 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA4 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA5 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA6 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA7 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA8 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA9 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA10 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA11 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA14 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOA15 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB4 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB5 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB6 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB7 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB8 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB9 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB10 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB11 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB13 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB14 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/DOB15 ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/RSTANOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/RSTBNOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/WEANOT ;
    wire \bridge/pci_target_unit/fifos/dpram16_3/INT_SIG ;
    wire \AD[27]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[26]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[25]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[24]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[23]/OUTBUF_GTS_AND_1_INV ;
    wire \CBE[3]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[17]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[16]/OUTBUF_GTS_AND_1_INV ;
    wire \CBE[2]/OUTBUF_GTS_AND_1_INV ;
    wire \STOP/OUTBUF_GTS_AND_1_INV ;
    wire \AD[22]/OUTBUF_GTS_AND_1_INV ;
    wire \FRAME/OUTBUF_GTS_AND_1_INV ;
    wire \PERR/OUTBUF_GTS_AND_1_INV ;
    wire \AD[21]/OUTBUF_GTS_AND_1_INV ;
    wire \IRDY/OUTBUF_GTS_AND_1_INV ;
    wire \AD[20]/OUTBUF_GTS_AND_1_INV ;
    wire \SERR/OUTBUF_GTS_AND_1_INV ;
    wire \AD[19]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[13]/OUTBUF_GTS_AND_1_INV ;
    wire \PAR/OUTBUF_GTS_AND_1_INV ;
    wire \AD[18]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[12]/OUTBUF_GTS_AND_1_INV ;
    wire \CBE[1]/OUTBUF_GTS_AND_1_INV ;
    wire \TRDY/OUTBUF_GTS_AND_1_INV ;
    wire \AD[11]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[15]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[14]/OUTBUF_GTS_AND_1_INV ;
    wire \DEVSEL/OUTBUF_GTS_AND_1_INV ;
    wire \AD[10]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[3]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[9]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[2]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[8]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[1]/OUTBUF_GTS_AND_1_INV ;
    wire \CBE[0]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[6]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[7]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[5]/OUTBUF_GTS_AND_1_INV ;
    wire C_HSYNC_2_INV;
    wire \AD[4]/OUTBUF_GTS_AND_1_INV ;
    wire \REQ/OUTBUF_GTS_AND_1_INV ;
    wire \AD[0]/OUTBUF_GTS_AND_1_INV ;
    wire C_VSYNC_2_INV;
    wire C_LED_2_INV;
    wire \AD[31]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[30]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[29]/OUTBUF_GTS_AND_1_INV ;
    wire \AD[28]/OUTBUF_GTS_AND_1_INV ;
    wire \C_RGB[14]_2_INV ;
    wire \C_RGB[7]_2_INV ;
    wire \C_RGB[15]_2_INV ;
    wire \C_RGB[8]_2_INV ;
    wire \C_RGB[9]_2_INV ;
    wire \C_RGB[4]_2_INV ;
    wire \C_RGB[5]_2_INV ;
    wire \C_RGB[10]_2_INV ;
    wire \C_RGB[6]_2_INV ;
    wire \C_RGB[11]_2_INV ;
    wire \C_RGB[12]_2_INV ;
    wire \C_RGB[13]_2_INV ;
    wire GND;
    wire VCC;
    wire GSR = glbl.GSR;
    wire GTS = glbl.GTS;
    wire [31:0] \bridge/pci_target_unit/pci_target_if/address1_in ;
    wire [31:0] \bridge/out_bckp_ad_out ;
    wire [31:0] \bridge/wishbone_slave_unit/pcim_if_address_out ;
    wire [31:2] \bridge/wishbone_slave_unit/wb_addr_dec/addr1 ;
    wire [31:2] \bridge/wishbone_slave_unit/wbs_sm_data_out ;
    wire [31:2] \bridge/wishbone_slave_unit/del_sync_addr_out ;
    wire [7:0] \bridge/pci_target_unit/wishbone_master/rty_counter ;
    wire [31:0] \bridge/pci_target_unit/fifos_pcir_data_out ;
    wire [31:0] \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg ;
    wire [31:0] \bridge/pci_target_unit/fifos_pciw_addr_data_out ;
    wire [31:0] \bridge/pci_target_unit/del_sync_addr_out ;
    wire [10:2] ADR_O;
    wire [3:2] \bridge/wishbone_slave_unit/wbs_sm_cbe_out ;
    wire [2:0] \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next ;
    wire [7:0] \bridge/conf_latency_tim_out ;
    wire [7:0] \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_raddr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_raddr_0 ;
    wire [5:0] \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr ;
    wire [5:0] \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one ;
    wire [5:0] \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one ;
    wire [3:0] \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 ;
    wire [2:0] \bridge/pci_target_unit/fifos/inNextGreyCount ;
    wire [3:0] \bridge/pci_target_unit/fifos/pciw_inTransactionCount ;
    wire [3:0] \bridge/pci_target_unit/fifos/inGreyCount ;
    wire [0:0] \bridge/conf_pci_img_ctrl1_out ;
    wire [8:2] \bridge/pciu_conf_offset_out ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next ;
    wire [31:0] \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out ;
    wire [31:0] \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data ;
    wire [16:0] \bridge/pci_target_unit/del_sync/comp_cycle_count ;
    wire [16:0] \bridge/wishbone_slave_unit/del_sync/comp_cycle_count ;
    wire [31:0] \bridge/wishbone_slave_unit/fifos_wbr_data_out ;
    wire [2:0] \bridge/pci_target_unit/wishbone_master/c_state ;
    wire [3:0] \bridge/pci_target_unit/fifos_pciw_cbe_out ;
    wire [3:0] \bridge/pci_target_unit/del_sync_be_out ;
    wire [31:24] \bridge/configuration/pci_err_cs_bit31_24 ;
    wire [3:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_waddr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next ;
    wire [3:0] \bridge/wishbone_slave_unit/pcim_if_be_out ;
    wire [3:0] \bridge/wishbone_slave_unit/pcim_if_next_be_out ;
    wire [3:0] \bridge/wishbone_slave_unit/pcim_if_bc_out ;
    wire [3:0] \bridge/pci_mux_cbe_in ;
    wire [3:0] \bridge/out_bckp_cbe_out ;
    wire [1:0] \bridge/pci_target_unit/fifos_pcir_control_out ;
    wire [1:0] \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg ;
    wire [1:0] \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out ;
    wire [3:0] \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt ;
    wire [9:0] \CRT/ssvga_fifo/rd_ptr_plus1 ;
    wire [9:0] \CRT/ssvga_fifo/rd_ptr ;
    wire [31:2] \CRT/pix_start_addr ;
    wire [1:0] \bridge/wishbone_slave_unit/pcim_if_wbr_control_out ;
    wire [3:1] \bridge/wishbone_slave_unit/del_sync_bc_out ;
    wire [3:0] \bridge/wishbone_slave_unit/fifos_wbw_cbe_out ;
    wire [0:0] \bridge/wishbone_slave_unit/wishbone_slave/img_hit ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_waddr ;
    wire [3:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbw_waddr ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next ;
    wire [3:0] \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be ;
    wire [3:0] \bridge/pci_target_unit/del_sync_bc_out ;
    wire [2:0] \bridge/wishbone_slave_unit/fifos/inNextGreyCount ;
    wire [3:0] \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount ;
    wire [3:0] \bridge/wishbone_slave_unit/fifos/inGreyCount ;
    wire [16:0] \CRT/ssvga_wbm_if/vmaddr_r ;
    wire [1:0] \bridge/pci_target_unit/pci_target_sm/c_state ;
    wire [0:0] \bridge/wishbone_slave_unit/fifos_wbw_control_out ;
    wire [3:3] \bridge/wishbone_slave_unit/wbs_sm_del_bc_out ;
    wire [3:0] \bridge/pci_target_unit/fifos/outGreyCount ;
    wire [0:0] \bridge/pci_target_unit/fifos_pciw_control_out ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 ;
    wire [9:0] \CRT/ssvga_crtc/hcntr ;
    wire [3:0] \bridge/wishbone_slave_unit/pcim_if_wbr_be_out ;
    wire [3:0] N_CBE;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr ;
    wire [5:0] \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr ;
    wire [5:0] \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr ;
    wire [3:0] \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 ;
    wire [9:0] \CRT/ssvga_crtc/vcntr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 ;
    wire [2:0] \bridge/pci_target_unit/fifos/outNextGreyCount ;
    wire [3:0] \bridge/pci_target_unit/fifos/pciw_outTransactionCount ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_raddr ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_raddr_0 ;
    wire [31:0] \bridge/wishbone_slave_unit/pcim_sm_data_out ;
    wire [9:9] \bridge/configuration/wb_err_cs_bit10_8 ;
    wire [1:0] \bridge/wishbone_slave_unit/fifos_wbr_control_out ;
    wire [2:0] \bridge/wishbone_slave_unit/wishbone_slave/c_state ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next ;
    wire [5:0] \bridge/wishbone_slave_unit/fifos/wbr_waddr ;
    wire [5:0] \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next ;
    wire [19:12] \bridge/conf_pci_ba0_out ;
    wire [9:0] \CRT/ssvga_fifo/sync_gray_rd_ptr ;
    wire [7:0] \bridge/conf_cache_line_size_out ;
    wire [8:0] \bridge/wishbone_slave_unit/pci_initiator_if/read_count ;
    wire [31:0] \bridge/wishbone_slave_unit/pcim_if_next_data_out ;
    wire [31:0] \bridge/wishbone_slave_unit/pcim_if_data_out ;
    wire [7:0] \CRT/ssvga_fifo/wr_ptr_plus1 ;
    wire [7:0] \CRT/ssvga_fifo/wr_ptr ;
    wire [3:0] \bridge/in_reg_cbe_out ;
    wire [19:12] \bridge/conf_pci_ba1_out ;
    wire [19:12] \bridge/conf_pci_am1_out ;
    wire [15:11] \bridge/configuration/status_bit15_11 ;
    wire [31:0] SDAT_O;
    wire [31:12] \bridge/configuration/pci_tran_addr1 ;
    wire [31:24] \bridge/configuration/wb_err_cs_bit31_24 ;
    wire [31:0] \bridge/configuration/pci_err_addr ;
    wire [19:12] \bridge/conf_wb_ba1_out ;
    wire [19:12] \bridge/conf_wb_am1_out ;
    wire [31:12] \bridge/configuration/wb_tran_addr1 ;
    wire [31:0] \bridge/configuration/pci_err_data ;
    wire [31:0] \bridge/configuration/wb_err_data ;
    wire [31:0] \bridge/configuration/wb_err_addr ;
    wire [23:12] \bridge/configuration/pci_addr_mask1 ;
    wire [23:12] \bridge/configuration/wb_base_addr1 ;
    wire [23:12] \bridge/configuration/wb_addr_mask1 ;
    wire [23:12] \bridge/configuration/pci_base_addr1 ;
    wire [23:12] \bridge/configuration/pci_base_addr0 ;
    wire [7:0] \bridge/configuration/interrupt_line ;
    wire [1:1] \bridge/conf_wb_img_ctrl1_out ;
    wire [9:0] \CRT/ssvga_fifo/gray_read_ptr ;
    wire [1:0] \bridge/pci_target_unit/pci_target_if/conf_addr_out ;
    wire [7:0] \bridge/pci_target_unit/wishbone_master/cache_line ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next ;
    wire [3:0] \bridge/pciu_err_bc_out ;
    wire [31:0] \bridge/pci_target_unit/pcit_if_addr_out ;
    wire [2:2] \bridge/configuration/pci_img_ctrl1 ;
    wire [4:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 ;
    wire [4:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 ;
    wire [3:0] \bridge/pci_target_unit/pcit_if_bc_out ;
    wire [7:0] \CRT/ssvga_fifo/dat_o_high ;
    wire [7:0] \CRT/ssvga_fifo/dat_o_low ;
    wire [7:0] \CRT/fifo_out ;
    wire [3:0] \bridge/wishbone_slave_unit/fifos/outGreyCount ;
    wire [31:0] \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out ;
    wire [3:0] \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out ;
    wire [15:4] \CRT/pal_pix_dat ;
    wire [15:4] rgb_int;
    wire [15:0] \CRT/wbs_pal_data ;
    wire [31:0] \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out ;
    wire [0:0] \bridge/wishbone_slave_unit/wbs_sm_wbw_control_out ;
    wire [3:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next ;
    wire [2:0] \bridge/wishbone_slave_unit/fifos/outNextGreyCount ;
    wire [4:0] \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next ;
    wire [3:0] \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next ;
    wire [3:0] \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next ;
    wire [1:1] \bridge/wishbone_slave_unit/amux_hit_out ;
    wire [3:0] \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next ;
    wire [8:0] \CRT/ssvga_fifo/gray_rd_ptr ;
    wire [31:0] N_AD;
    wire [31:0] AD_out;
    wire [31:0] AD_en;
    wire [3:0] CBE_out;
    wire [3:0] CBE_en;
    wire [15:4] N_RGB;
    initial $sdf_annotate("crt_time_sim.sdf");
    defparam C18859.INIT = 16'hA0A0;
    X_LUT4 C18859(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .ADR3 (VCC),
      .O (\bridge/configuration/delete_pci_err_cs_bit10/GROM )
    );
    defparam C18831.INIT = 16'h8888;
    X_LUT4 C18831(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [10]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/configuration/C387/N3 )
    );
    X_INV \bridge/configuration/delete_pci_err_cs_bit10/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/delete_pci_err_cs_bit10/SRNOT )
    );
    X_BUF \bridge/configuration/delete_pci_err_cs_bit10/YUSED (
      .I (\bridge/configuration/delete_pci_err_cs_bit10/GROM ),
      .O (\bridge/configuration/C390/N3 )
    );
    X_FF \bridge/configuration/delete_pci_err_cs_bit8_reg (
      .I (\bridge/configuration/delete_pci_err_cs_bit10/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C343/N5 ),
      .SET (\bridge/configuration/delete_pci_err_cs_bit10/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_pci_err_cs_bit8 )
    );
    X_OR2 \bridge/configuration/delete_pci_err_cs_bit10/FFY/ASYNC_FF_GSR_OR_0 (
      .I0 (\bridge/configuration/delete_pci_err_cs_bit10/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_pci_err_cs_bit10/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/delete_pci_err_cs_bit10_reg (
      .I (\bridge/configuration/C387/N3 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C343/N5 ),
      .SET (\bridge/configuration/delete_pci_err_cs_bit10/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_pci_err_cs_bit10 )
    );
    X_OR2 \bridge/configuration/delete_pci_err_cs_bit10/FFX/ASYNC_FF_GSR_OR_1 (
      .I0 (\bridge/configuration/delete_pci_err_cs_bit10/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_pci_err_cs_bit10/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18761.INIT = 16'hFFFE;
    X_LUT4 C18761(
      .ADR0 (syn20486),
      .ADR1 (syn20502),
      .ADR2 (syn179882),
      .ADR3 (syn179883),
      .O (\bridge/out_bckp_ad_out[0]/GROM )
    );
    defparam C18762.INIT = 16'hFEEE;
    X_LUT4 C18762(
      .ADR0 (syn179881),
      .ADR1 (syn179878),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn17116),
      .O (\bridge/out_bckp_ad_out[0]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[0]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<0>/YUSED (
      .I (\bridge/out_bckp_ad_out[0]/GROM ),
      .O (\bridge/output_backup/C3/N6 )
    );
    X_BUF \bridge/out_bckp_ad_out<0>/XUSED (
      .I (\bridge/out_bckp_ad_out[0]/FROM ),
      .O (syn179883)
    );
    X_FF \bridge/output_backup/ad_out_reg<0> (
      .I (\bridge/out_bckp_ad_out[0]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [0])
    );
    X_OR2 \bridge/out_bckp_ad_out<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18747.INIT = 16'hBB88;
    X_LUT4 C18747(
      .ADR0 (syn20532),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (VCC),
      .ADR3 (syn20538),
      .O (\bridge/out_bckp_ad_out[1]/GROM )
    );
    defparam C18748.INIT = 16'hECEC;
    X_LUT4 C18748(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [1]),
      .ADR1 (syn179894),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR3 (VCC),
      .O (\bridge/out_bckp_ad_out[1]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[1]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<1>/YUSED (
      .I (\bridge/out_bckp_ad_out[1]/GROM ),
      .O (\bridge/output_backup/C3/N12 )
    );
    X_BUF \bridge/out_bckp_ad_out<1>/XUSED (
      .I (\bridge/out_bckp_ad_out[1]/FROM ),
      .O (syn20538)
    );
    X_FF \bridge/output_backup/ad_out_reg<1> (
      .I (\bridge/out_bckp_ad_out[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [1])
    );
    X_OR2 \bridge/out_bckp_ad_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19347.INIT = 16'h8000;
    X_LUT4 C19347(
      .ADR0 (syn177396),
      .ADR1 (N12360),
      .ADR2 (syn177397),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/GROM )
    );
    defparam C19348.INIT = 16'h8000;
    X_LUT4 C19348(
      .ADR0 (syn177396),
      .ADR1 (N12360),
      .ADR2 (syn177397),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<3>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [2])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<3>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [3])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<2> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [2])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_addr_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<3> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [3])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_addr_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18734.INIT = 16'hEFE0;
    X_LUT4 C18734(
      .ADR0 (syn179960),
      .ADR1 (syn20564),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn20571),
      .O (\bridge/out_bckp_ad_out[2]/GROM )
    );
    defparam C18738.INIT = 16'hFCF0;
    X_LUT4 C18738(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [2]),
      .ADR2 (syn179931),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\bridge/out_bckp_ad_out[2]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[2]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<2>/YUSED (
      .I (\bridge/out_bckp_ad_out[2]/GROM ),
      .O (\bridge/output_backup/C3/N18 )
    );
    X_BUF \bridge/out_bckp_ad_out<2>/XUSED (
      .I (\bridge/out_bckp_ad_out[2]/FROM ),
      .O (syn20571)
    );
    X_FF \bridge/output_backup/ad_out_reg<2> (
      .I (\bridge/out_bckp_ad_out[2]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[2]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [2])
    );
    X_OR2 \bridge/out_bckp_ad_out<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[2]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17814.INIT = 16'h0F0C;
    X_LUT4 C17814(
      .ADR0 (VCC),
      .ADR1 (syn19555),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3068 ),
      .O (\bridge/pci_target_unit/wishbone_master/C107/N5 )
    );
    defparam C17811.INIT = 16'h5544;
    X_LUT4 C17811(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .ADR1 (syn19555),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3069 ),
      .O (\bridge/pci_target_unit/wishbone_master/C107/N10 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/rty_counter<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/rty_counter_reg<0> (
      .I (\bridge/pci_target_unit/wishbone_master/C107/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter [0])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/rty_counter<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/rty_counter[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/rty_counter_reg<1> (
      .I (\bridge/pci_target_unit/wishbone_master/C107/N10 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter [1])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/rty_counter<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/rty_counter[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18715.INIT = 16'hFEEE;
    X_LUT4 C18715(
      .ADR0 (syn20611),
      .ADR1 (syn180003),
      .ADR2 (syn20598),
      .ADR3 (syn180250),
      .O (\bridge/out_bckp_ad_out[3]/GROM )
    );
    defparam C18716.INIT = 16'hA0A0;
    X_LUT4 C18716(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (VCC),
      .ADR2 (syn17106),
      .ADR3 (VCC),
      .O (\bridge/out_bckp_ad_out[3]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[3]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<3>/YUSED (
      .I (\bridge/out_bckp_ad_out[3]/GROM ),
      .O (\bridge/output_backup/C3/N24 )
    );
    X_BUF \bridge/out_bckp_ad_out<3>/XUSED (
      .I (\bridge/out_bckp_ad_out[3]/FROM ),
      .O (syn180250)
    );
    X_FF \bridge/output_backup/ad_out_reg<3> (
      .I (\bridge/out_bckp_ad_out[3]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [3])
    );
    X_OR2 \bridge/out_bckp_ad_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17782.INIT = 16'h0A0A;
    X_LUT4 C17782(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/norm_prf_en ),
      .ADR1 (VCC),
      .ADR2 (\bridge/in_reg_frame_out ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/pcit_if_burst_out )
    );
    defparam C19216.INIT = 16'hFCCC;
    X_LUT4 C19216(
      .ADR0 (VCC),
      .ADR1 (syn19671),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR3 (\bridge/in_reg_frame_out ),
      .O (\bridge/pci_target_unit/del_sync_burst_out/FROM )
    );
    X_INV \bridge/pci_target_unit/del_sync_burst_out/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_burst_out/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/del_sync_burst_out/XUSED (
      .I (\bridge/pci_target_unit/del_sync_burst_out/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_control_out[0] )
    );
    X_FF \bridge/pci_target_unit/del_sync/burst_out_reg (
      .I (\bridge/pci_target_unit/pcit_if_burst_out ),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_burst_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_burst_out )
    );
    X_OR2 \bridge/pci_target_unit/del_sync_burst_out/FFY/ASYNC_FF_GSR_OR_2 (
      .I0 (\bridge/pci_target_unit/del_sync_burst_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_burst_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19349.INIT = 16'h8000;
    X_LUT4 C19349(
      .ADR0 (syn177396),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR2 (syn177397),
      .ADR3 (N12360),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/GROM )
    );
    defparam C19350.INIT = 16'h8080;
    X_LUT4 C19350(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR2 (N12360),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<5>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [4])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<5>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [5])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<4> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [4])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_addr_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<5> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [5])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_addr_out<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18701.INIT = 16'hAFA0;
    X_LUT4 C18701(
      .ADR0 (syn20635),
      .ADR1 (VCC),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn20641),
      .O (\bridge/out_bckp_ad_out[4]/GROM )
    );
    defparam C18702.INIT = 16'hFAAA;
    X_LUT4 C18702(
      .ADR0 (syn180012),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [4]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\bridge/out_bckp_ad_out[4]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[4]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<4>/YUSED (
      .I (\bridge/out_bckp_ad_out[4]/GROM ),
      .O (\bridge/output_backup/C3/N30 )
    );
    X_BUF \bridge/out_bckp_ad_out<4>/XUSED (
      .I (\bridge/out_bckp_ad_out[4]/FROM ),
      .O (syn20641)
    );
    X_FF \bridge/output_backup/ad_out_reg<4> (
      .I (\bridge/out_bckp_ad_out[4]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [4])
    );
    X_OR2 \bridge/out_bckp_ad_out<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[4]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17810.INIT = 16'h5550;
    X_LUT4 C17810(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/N3070 ),
      .ADR3 (syn19555),
      .O (\bridge/pci_target_unit/wishbone_master/C107/N15 )
    );
    defparam C17809.INIT = 16'h00EE;
    X_LUT4 C17809(
      .ADR0 (syn19555),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3071 ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .O (\bridge/pci_target_unit/wishbone_master/C107/N20 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/rty_counter<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/rty_counter_reg<2> (
      .I (\bridge/pci_target_unit/wishbone_master/C107/N15 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter [2])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/rty_counter<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/rty_counter[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/rty_counter_reg<3> (
      .I (\bridge/pci_target_unit/wishbone_master/C107/N20 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter [3])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/rty_counter<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/rty_counter[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18689.INIT = 16'hFFFA;
    X_LUT4 C18689(
      .ADR0 (syn20662),
      .ADR1 (VCC),
      .ADR2 (syn20672),
      .ADR3 (syn180067),
      .O (\bridge/out_bckp_ad_out[5]/GROM )
    );
    defparam C18690.INIT = 16'hEAC0;
    X_LUT4 C18690(
      .ADR0 (syn136386),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [5]),
      .ADR2 (syn136384),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [5]),
      .O (\bridge/out_bckp_ad_out[5]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[5]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<5>/YUSED (
      .I (\bridge/out_bckp_ad_out[5]/GROM ),
      .O (\bridge/output_backup/C3/N36 )
    );
    X_BUF \bridge/out_bckp_ad_out<5>/XUSED (
      .I (\bridge/out_bckp_ad_out[5]/FROM ),
      .O (syn180067)
    );
    X_FF \bridge/output_backup/ad_out_reg<5> (
      .I (\bridge/out_bckp_ad_out[5]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [5])
    );
    X_OR2 \bridge/out_bckp_ad_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19352.INIT = 16'h8000;
    X_LUT4 C19352(
      .ADR0 (N12360),
      .ADR1 (syn177397),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR3 (syn177396),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/GROM )
    );
    defparam C19353.INIT = 16'h8000;
    X_LUT4 C19353(
      .ADR0 (syn177396),
      .ADR1 (syn177397),
      .ADR2 (N12360),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<7>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [6])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<7>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [7])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<6> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [6])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_addr_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<7> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [7])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_addr_out<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18679.INIT = 16'hFFEA;
    X_LUT4 C18679(
      .ADR0 (syn180098),
      .ADR1 (syn20688),
      .ADR2 (syn180250),
      .ADR3 (syn20701),
      .O (\bridge/out_bckp_ad_out[6]/GROM )
    );
    X_INV \bridge/out_bckp_ad_out<6>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[6]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<6>/YUSED (
      .I (\bridge/out_bckp_ad_out[6]/GROM ),
      .O (\bridge/output_backup/C3/N42 )
    );
    X_FF \bridge/output_backup/ad_out_reg<6> (
      .I (\bridge/out_bckp_ad_out[6]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[6]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [6])
    );
    X_OR2 \bridge/out_bckp_ad_out<6>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[6]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[6]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17808.INIT = 16'h0F0A;
    X_LUT4 C17808(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3072 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .ADR3 (syn19555),
      .O (\bridge/pci_target_unit/wishbone_master/C107/N25 )
    );
    defparam C17807.INIT = 16'h0F0C;
    X_LUT4 C17807(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3073 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .ADR3 (syn19555),
      .O (\bridge/pci_target_unit/wishbone_master/C107/N30 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/rty_counter<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter[5]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/rty_counter_reg<4> (
      .I (\bridge/pci_target_unit/wishbone_master/C107/N25 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter [4])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/rty_counter<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/rty_counter[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/rty_counter_reg<5> (
      .I (\bridge/pci_target_unit/wishbone_master/C107/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter [5])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/rty_counter<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/rty_counter[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17869.INIT = 16'hFF88;
    X_LUT4 C17869(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [10]),
      .ADR1 (syn16925),
      .ADR2 (VCC),
      .ADR3 (syn182174),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N66 )
    );
    defparam C17870.INIT = 16'hB3A0;
    X_LUT4 C17870(
      .ADR0 (syn16933),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [10]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N2993 ),
      .O (\ADR_O[10]/FROM )
    );
    X_INV \ADR_O<10>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[10]/SRNOT )
    );
    X_BUF \ADR_O<10>/XUSED (
      .I (\ADR_O[10]/FROM ),
      .O (syn182174)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<10> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N66 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[10]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[10])
    );
    X_OR2 \ADR_O<10>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[10]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[10]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18669.INIT = 16'hCFC0;
    X_LUT4 C18669(
      .ADR0 (VCC),
      .ADR1 (syn20720),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn20726),
      .O (\bridge/out_bckp_ad_out[7]/GROM )
    );
    defparam C18670.INIT = 16'hFAF0;
    X_LUT4 C18670(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (VCC),
      .ADR2 (syn180107),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [7]),
      .O (\bridge/out_bckp_ad_out[7]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[7]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<7>/YUSED (
      .I (\bridge/out_bckp_ad_out[7]/GROM ),
      .O (\bridge/output_backup/C3/N48 )
    );
    X_BUF \bridge/out_bckp_ad_out<7>/XUSED (
      .I (\bridge/out_bckp_ad_out[7]/FROM ),
      .O (syn20726)
    );
    X_FF \bridge/output_backup/ad_out_reg<7> (
      .I (\bridge/out_bckp_ad_out[7]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [7])
    );
    X_OR2 \bridge/out_bckp_ad_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19354.INIT = 16'hF000;
    X_LUT4 C19354(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (N12360),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/GROM )
    );
    defparam C19670.INIT = 16'h8800;
    X_LUT4 C19670(
      .ADR0 (syn177396),
      .ADR1 (syn177397),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [8]),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<8>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<8>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [8])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<8>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/FROM ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<8> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [8])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_addr_out<8>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[8]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17867.INIT = 16'hFF88;
    X_LUT4 C17867(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [11]),
      .ADR1 (syn16925),
      .ADR2 (VCC),
      .ADR3 (syn182179),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N72 )
    );
    defparam C17868.INIT = 16'hAE0C;
    X_LUT4 C17868(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [11]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N2994 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR3 (syn16933),
      .O (\bridge/pciu_err_addr_out[11]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[11]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<11>/XUSED (
      .I (\bridge/pciu_err_addr_out[11]/FROM ),
      .O (syn182179)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<11> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N72 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[11] )
    );
    X_OR2 \bridge/pciu_err_addr_out<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[11]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18649.INIT = 16'hFFFE;
    X_LUT4 C18649(
      .ADR0 (syn20759),
      .ADR1 (syn180180),
      .ADR2 (syn180181),
      .ADR3 (syn180185),
      .O (\bridge/out_bckp_ad_out[8]/GROM )
    );
    defparam C18650.INIT = 16'hFFFE;
    X_LUT4 C18650(
      .ADR0 (syn180183),
      .ADR1 (syn20738),
      .ADR2 (syn20737),
      .ADR3 (syn180176),
      .O (\bridge/out_bckp_ad_out[8]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<8>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[8]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<8>/YUSED (
      .I (\bridge/out_bckp_ad_out[8]/GROM ),
      .O (\bridge/output_backup/C3/N54 )
    );
    X_BUF \bridge/out_bckp_ad_out<8>/XUSED (
      .I (\bridge/out_bckp_ad_out[8]/FROM ),
      .O (syn180185)
    );
    X_FF \bridge/output_backup/ad_out_reg<8> (
      .I (\bridge/out_bckp_ad_out[8]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[8]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [8])
    );
    X_OR2 \bridge/out_bckp_ad_out<8>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[8]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[8]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17806.INIT = 16'h0F0A;
    X_LUT4 C17806(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3074 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .ADR3 (syn19555),
      .O (\bridge/pci_target_unit/wishbone_master/C107/N35 )
    );
    defparam C17805.INIT = 16'h0E0E;
    X_LUT4 C17805(
      .ADR0 (syn19555),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3075 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/C107/N40 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/rty_counter<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter[7]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/rty_counter_reg<6> (
      .I (\bridge/pci_target_unit/wishbone_master/C107/N35 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter [6])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/rty_counter<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/rty_counter[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/rty_counter_reg<7> (
      .I (\bridge/pci_target_unit/wishbone_master/C107/N40 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_counter [7])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/rty_counter<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/rty_counter[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/rty_counter[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19355.INIT = 16'h8080;
    X_LUT4 C19355(
      .ADR0 (N12360),
      .ADR1 (syn24500),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [9]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/GROM )
    );
    defparam C19366.INIT = 16'h5F5F;
    X_LUT4 C19366(
      .ADR0 (N12360),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/map ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<9>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [9])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<9>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_cbe_out [2])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<9> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [9])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_addr_out<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[9]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17849.INIT = 16'hFFC0;
    X_LUT4 C17849(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [20]),
      .ADR2 (syn16925),
      .ADR3 (syn182224),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N126 )
    );
    defparam C17850.INIT = 16'hAE0C;
    X_LUT4 C17850(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [20]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3003 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR3 (syn16933),
      .O (\bridge/pciu_err_addr_out[20]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<20>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[20]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<20>/XUSED (
      .I (\bridge/pciu_err_addr_out[20]/FROM ),
      .O (syn182224)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<20> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N126 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[20]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[20] )
    );
    X_OR2 \bridge/pciu_err_addr_out<20>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[20]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[20]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17865.INIT = 16'hFFC0;
    X_LUT4 C17865(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [12]),
      .ADR2 (syn16925),
      .ADR3 (syn182184),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N78 )
    );
    defparam C17866.INIT = 16'hC0EA;
    X_LUT4 C17866(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N2995 ),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [12]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\bridge/pciu_err_addr_out[12]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<12>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[12]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<12>/XUSED (
      .I (\bridge/pciu_err_addr_out[12]/FROM ),
      .O (syn182184)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<12> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N78 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[12]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[12] )
    );
    X_OR2 \bridge/pciu_err_addr_out<12>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[12]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[12]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18633.INIT = 16'hFFEA;
    X_LUT4 C18633(
      .ADR0 (syn180222),
      .ADR1 (syn137911),
      .ADR2 (syn180212),
      .ADR3 (syn20788),
      .O (\bridge/out_bckp_ad_out[9]/GROM )
    );
    defparam C18646.INIT = 16'h00EC;
    X_LUT4 C18646(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (syn180219),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [9]),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\bridge/out_bckp_ad_out[9]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[9]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<9>/YUSED (
      .I (\bridge/out_bckp_ad_out[9]/GROM ),
      .O (\bridge/output_backup/C3/N60 )
    );
    X_BUF \bridge/out_bckp_ad_out<9>/XUSED (
      .I (\bridge/out_bckp_ad_out[9]/FROM ),
      .O (syn20788)
    );
    X_FF \bridge/output_backup/ad_out_reg<9> (
      .I (\bridge/out_bckp_ad_out[9]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [9])
    );
    X_OR2 \bridge/out_bckp_ad_out<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[9]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17847.INIT = 16'hFF88;
    X_LUT4 C17847(
      .ADR0 (syn16925),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [21]),
      .ADR2 (VCC),
      .ADR3 (syn182229),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N132 )
    );
    defparam C17848.INIT = 16'hF222;
    X_LUT4 C17848(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3004 ),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [21]),
      .ADR3 (syn16933),
      .O (\bridge/pciu_err_addr_out[21]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[21]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<21>/XUSED (
      .I (\bridge/pciu_err_addr_out[21]/FROM ),
      .O (syn182229)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<21> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N132 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[21] )
    );
    X_OR2 \bridge/pciu_err_addr_out<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[21]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17863.INIT = 16'hFFC0;
    X_LUT4 C17863(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [13]),
      .ADR2 (syn16925),
      .ADR3 (syn182189),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N84 )
    );
    defparam C17864.INIT = 16'hF444;
    X_LUT4 C17864(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N2996 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [13]),
      .ADR3 (syn16933),
      .O (\bridge/pciu_err_addr_out[13]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[13]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<13>/XUSED (
      .I (\bridge/pciu_err_addr_out[13]/FROM ),
      .O (syn182189)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<13> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N84 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[13] )
    );
    X_OR2 \bridge/pciu_err_addr_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17829.INIT = 16'hFFC0;
    X_LUT4 C17829(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [30]),
      .ADR2 (syn16925),
      .ADR3 (syn182274),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N186 )
    );
    defparam C17830.INIT = 16'hA0EC;
    X_LUT4 C17830(
      .ADR0 (syn16933),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3013 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [30]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\bridge/pciu_err_addr_out[30]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<30>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[30]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<30>/XUSED (
      .I (\bridge/pciu_err_addr_out[30]/FROM ),
      .O (syn182274)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<30> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N186 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[30]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[30] )
    );
    X_OR2 \bridge/pciu_err_addr_out<30>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[30]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[30]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17845.INIT = 16'hFF88;
    X_LUT4 C17845(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [22]),
      .ADR1 (syn16925),
      .ADR2 (VCC),
      .ADR3 (syn182234),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N138 )
    );
    defparam C17846.INIT = 16'h88F8;
    X_LUT4 C17846(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [22]),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/N3005 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\bridge/pciu_err_addr_out[22]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<22>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[22]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<22>/XUSED (
      .I (\bridge/pciu_err_addr_out[22]/FROM ),
      .O (syn182234)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<22> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N138 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[22]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[22] )
    );
    X_OR2 \bridge/pciu_err_addr_out<22>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[22]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[22]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17861.INIT = 16'hFF88;
    X_LUT4 C17861(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [14]),
      .ADR1 (syn16925),
      .ADR2 (VCC),
      .ADR3 (syn182194),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N90 )
    );
    defparam C17862.INIT = 16'h8F88;
    X_LUT4 C17862(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [14]),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N2997 ),
      .O (\bridge/pciu_err_addr_out[14]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<14>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[14]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<14>/XUSED (
      .I (\bridge/pciu_err_addr_out[14]/FROM ),
      .O (syn182194)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<14> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N90 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[14]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[14] )
    );
    X_OR2 \bridge/pciu_err_addr_out<14>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[14]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[14]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17827.INIT = 16'hFFC0;
    X_LUT4 C17827(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [31]),
      .ADR2 (syn16925),
      .ADR3 (syn182279),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N192 )
    );
    defparam C17828.INIT = 16'hF444;
    X_LUT4 C17828(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3014 ),
      .ADR2 (syn16933),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [31]),
      .O (\bridge/pciu_err_addr_out[31]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[31]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<31>/XUSED (
      .I (\bridge/pciu_err_addr_out[31]/FROM ),
      .O (syn182279)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<31> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N192 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[31] )
    );
    X_OR2 \bridge/pciu_err_addr_out<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[31]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17843.INIT = 16'hFFC0;
    X_LUT4 C17843(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [23]),
      .ADR2 (syn16925),
      .ADR3 (syn182239),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N144 )
    );
    defparam C17844.INIT = 16'hA0EC;
    X_LUT4 C17844(
      .ADR0 (syn16933),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3006 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [23]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\bridge/pciu_err_addr_out[23]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[23]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<23>/XUSED (
      .I (\bridge/pciu_err_addr_out[23]/FROM ),
      .O (syn182239)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<23> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N144 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[23] )
    );
    X_OR2 \bridge/pciu_err_addr_out<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[23]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17859.INIT = 16'hFFA0;
    X_LUT4 C17859(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [15]),
      .ADR1 (VCC),
      .ADR2 (syn16925),
      .ADR3 (syn182199),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N96 )
    );
    defparam C17860.INIT = 16'hA0EC;
    X_LUT4 C17860(
      .ADR0 (syn16933),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N2998 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [15]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\bridge/pciu_err_addr_out[15]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[15]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<15>/XUSED (
      .I (\bridge/pciu_err_addr_out[15]/FROM ),
      .O (syn182199)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<15> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N96 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[15] )
    );
    X_OR2 \bridge/pciu_err_addr_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17841.INIT = 16'hFFC0;
    X_LUT4 C17841(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [24]),
      .ADR2 (syn16925),
      .ADR3 (syn182244),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N150 )
    );
    defparam C17842.INIT = 16'hC0EA;
    X_LUT4 C17842(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3007 ),
      .ADR1 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [24]),
      .ADR2 (syn16933),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\bridge/pciu_err_addr_out[24]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<24>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[24]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<24>/XUSED (
      .I (\bridge/pciu_err_addr_out[24]/FROM ),
      .O (syn182244)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<24> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N150 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[24]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[24] )
    );
    X_OR2 \bridge/pciu_err_addr_out<24>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[24]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[24]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17857.INIT = 16'hFF88;
    X_LUT4 C17857(
      .ADR0 (syn16925),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [16]),
      .ADR2 (VCC),
      .ADR3 (syn182204),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N102 )
    );
    defparam C17858.INIT = 16'h88F8;
    X_LUT4 C17858(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [16]),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/N2999 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\bridge/pciu_err_addr_out[16]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<16>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[16]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<16>/XUSED (
      .I (\bridge/pciu_err_addr_out[16]/FROM ),
      .O (syn182204)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<16> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N102 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[16]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[16] )
    );
    X_OR2 \bridge/pciu_err_addr_out<16>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[16]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[16]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17839.INIT = 16'hFFC0;
    X_LUT4 C17839(
      .ADR0 (VCC),
      .ADR1 (syn16925),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [25]),
      .ADR3 (syn182249),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N156 )
    );
    defparam C17840.INIT = 16'hB3A0;
    X_LUT4 C17840(
      .ADR0 (syn16933),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [25]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3008 ),
      .O (\bridge/pciu_err_addr_out[25]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[25]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<25>/XUSED (
      .I (\bridge/pciu_err_addr_out[25]/FROM ),
      .O (syn182249)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<25> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N156 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[25] )
    );
    X_OR2 \bridge/pciu_err_addr_out<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[25]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17855.INIT = 16'hFFA0;
    X_LUT4 C17855(
      .ADR0 (syn16925),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [17]),
      .ADR3 (syn182209),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N108 )
    );
    defparam C17856.INIT = 16'hD5C0;
    X_LUT4 C17856(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [17]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3000 ),
      .O (\bridge/pciu_err_addr_out[17]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[17]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<17>/XUSED (
      .I (\bridge/pciu_err_addr_out[17]/FROM ),
      .O (syn182209)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<17> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N108 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[17] )
    );
    X_OR2 \bridge/pciu_err_addr_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17837.INIT = 16'hFF88;
    X_LUT4 C17837(
      .ADR0 (syn16925),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [26]),
      .ADR2 (VCC),
      .ADR3 (syn182254),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N162 )
    );
    defparam C17838.INIT = 16'hCE0A;
    X_LUT4 C17838(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3009 ),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [26]),
      .O (\bridge/pciu_err_addr_out[26]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<26>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[26]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<26>/XUSED (
      .I (\bridge/pciu_err_addr_out[26]/FROM ),
      .O (syn182254)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<26> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N162 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[26]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[26] )
    );
    X_OR2 \bridge/pciu_err_addr_out<26>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[26]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[26]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17853.INIT = 16'hFFA0;
    X_LUT4 C17853(
      .ADR0 (syn16925),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [18]),
      .ADR3 (syn182214),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N114 )
    );
    defparam C17854.INIT = 16'hA0EC;
    X_LUT4 C17854(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [18]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3001 ),
      .ADR2 (syn16933),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\bridge/pciu_err_addr_out[18]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<18>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[18]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<18>/XUSED (
      .I (\bridge/pciu_err_addr_out[18]/FROM ),
      .O (syn182214)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<18> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N114 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[18]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[18] )
    );
    X_OR2 \bridge/pciu_err_addr_out<18>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[18]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[18]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18220.INIT = 16'h3300;
    X_LUT4 C18220(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [0]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_13/cell0 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N5 )
    );
    defparam C18221.INIT = 16'h8000;
    X_LUT4 C18221(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (N_DEVSEL),
      .ADR2 (N_TRDY),
      .ADR3 (N_STOP),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/S_13/cell0 )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count_reg<0> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[0]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_stop_critical/C54 .INIT = 16'h04FF;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_stop_critical/C54 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/stop_w ),
      .ADR1 (N_IRDY),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/stop_w_frm ),
      .ADR3 
      (\bridge/pci_target_unit/pci_target_sm/pci_target_stop_critical/syn67 ),
      .O (\bridge/out_bckp_stop_out/GROM )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_stop_critical/C55 .INIT = 16'hFF54;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_stop_critical/C55 (
      .ADR0 (N_FRAME),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/stop_w_frm ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/stop_w ),
      .O (\bridge/out_bckp_stop_out/FROM )
    );
    X_INV \bridge/out_bckp_stop_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_stop_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_stop_out/YUSED (
      .I (\bridge/out_bckp_stop_out/GROM ),
      .O (N12476)
    );
    X_BUF \bridge/out_bckp_stop_out/XUSED (
      .I (\bridge/out_bckp_stop_out/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/pci_target_stop_critical/syn67 )
    );
    X_FF \bridge/output_backup/stop_out_reg (
      .I (\bridge/out_bckp_stop_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\bridge/out_bckp_stop_out/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_stop_out )
    );
    X_OR2 \bridge/out_bckp_stop_out/FFY/ASYNC_FF_GSR_OR_3 (
      .I0 (\bridge/out_bckp_stop_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_stop_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17835.INIT = 16'hFFC0;
    X_LUT4 C17835(
      .ADR0 (VCC),
      .ADR1 (syn16925),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [27]),
      .ADR3 (syn182259),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N168 )
    );
    defparam C17836.INIT = 16'hF222;
    X_LUT4 C17836(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3010 ),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR2 (syn16933),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [27]),
      .O (\bridge/pciu_err_addr_out[27]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[27]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<27>/XUSED (
      .I (\bridge/pciu_err_addr_out[27]/FROM ),
      .O (syn182259)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<27> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N168 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[27] )
    );
    X_OR2 \bridge/pciu_err_addr_out<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[27]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17851.INIT = 16'hFF88;
    X_LUT4 C17851(
      .ADR0 (syn16925),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [19]),
      .ADR2 (VCC),
      .ADR3 (syn182219),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N120 )
    );
    defparam C17852.INIT = 16'hBA30;
    X_LUT4 C17852(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [19]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/N3002 ),
      .ADR3 (syn16933),
      .O (\bridge/pciu_err_addr_out[19]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[19]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<19>/XUSED (
      .I (\bridge/pciu_err_addr_out[19]/FROM ),
      .O (syn182219)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<19> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N120 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[19] )
    );
    X_OR2 \bridge/pciu_err_addr_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18214.INIT = 16'hA00A;
    X_LUT4 C18214(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_13/cell0 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [0]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [1]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N10 )
    );
    defparam C18216.INIT = 16'hE1FF;
    X_LUT4 C18216(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [1]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [0]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [2]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_13/cell0 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N17 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count_reg<1> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N10 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count_reg<2> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2704/N17 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/decode_count<2>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count[2]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17833.INIT = 16'hFFC0;
    X_LUT4 C17833(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [28]),
      .ADR2 (syn16925),
      .ADR3 (syn182264),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N174 )
    );
    defparam C17834.INIT = 16'hB3A0;
    X_LUT4 C17834(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [28]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR2 (syn16933),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3011 ),
      .O (\bridge/pciu_err_addr_out[28]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<28>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[28]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<28>/XUSED (
      .I (\bridge/pciu_err_addr_out[28]/FROM ),
      .O (syn182264)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<28> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N174 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[28]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[28] )
    );
    X_OR2 \bridge/pciu_err_addr_out<28>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[28]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[28]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17628.INIT = 16'hFF0A;
    X_LUT4 C17628(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0 ),
      .ADR1 (VCC),
      .ADR2 (N12616),
      .ADR3 (syn23757),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_full )
    );
    defparam C17629.INIT = 16'h8200;
    X_LUT4 C17629(
      .ADR0 (syn182641),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [0]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [0]),
      .ADR3 (syn182642),
      .O (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FROM ),
      .O (syn23757)
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/full_reg (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_full ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos_pciw_full_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FFY/ASYNC_FF_GSR_OR_4 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FFX/ASYNC_FF_GSR_OR_5 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17831.INIT = 16'hFFA0;
    X_LUT4 C17831(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [29]),
      .ADR1 (VCC),
      .ADR2 (syn16925),
      .ADR3 (syn182269),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N180 )
    );
    defparam C17832.INIT = 16'hCE0A;
    X_LUT4 C17832(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3012 ),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [29]),
      .O (\bridge/pciu_err_addr_out[29]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[29]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<29>/XUSED (
      .I (\bridge/pciu_err_addr_out[29]/FROM ),
      .O (syn182269)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<29> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N180 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[29] )
    );
    X_OR2 \bridge/pciu_err_addr_out<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[29]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18213.INIT = 16'hF0AA;
    X_LUT4 C18213(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/conf_latency_tim_out [0]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N6 )
    );
    defparam C18211.INIT = 16'hF0CC;
    X_LUT4 C18211(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2619 ),
      .ADR2 (\bridge/conf_latency_tim_out [1]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N12 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer_reg<0> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12351),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer_reg<1> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (N12351),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19237.INIT = 16'hCCD8;
    X_LUT4 C19237(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [0]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [0]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/GROM )
    );
    defparam C19240.INIT = 16'hFE02;
    X_LUT4 C19240(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [1]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty ),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [1]),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_raddr_0<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_raddr_0<1>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/GROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr [0])
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_raddr_0<1>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr [1])
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_raddr_0_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0 [0])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_raddr_0<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_raddr_0_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0 [1])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_raddr_0<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18210.INIT = 16'hFA0A;
    X_LUT4 C18210(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2620 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .ADR3 (\bridge/conf_latency_tim_out [2]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N18 )
    );
    defparam C18209.INIT = 16'hE4E4;
    X_LUT4 C18209(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2621 ),
      .ADR2 (\bridge/conf_latency_tim_out [3]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N24 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer_reg<2> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (N12351),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer_reg<3> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N24 ),
      .CLK (CLK_BUFGPed),
      .CE (N12351),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19243.INIT = 16'hFE10;
    X_LUT4 C19243(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty ),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [2]),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/GROM )
    );
    defparam C19246.INIT = 16'hF0E2;
    X_LUT4 C19246(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_raddr_0<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_raddr_0<3>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/GROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr [2])
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_raddr_0<3>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr [3])
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_raddr_0_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0 [2])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_raddr_0<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_raddr_0_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0 [3])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_raddr_0<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18208.INIT = 16'hF0AA;
    X_LUT4 C18208(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2622 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/conf_latency_tim_out [4]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N30 )
    );
    defparam C18207.INIT = 16'hFC0C;
    X_LUT4 C18207(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2623 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .ADR3 (\bridge/conf_latency_tim_out [5]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N36 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer_reg<4> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (N12351),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer_reg<5> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (N12351),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [5])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[5]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19249.INIT = 16'hAAAC;
    X_LUT4 C19249(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[4]/GROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_raddr_0<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[4]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_raddr_0<4>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[4]/GROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr [4])
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_raddr_0_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_raddr_0[4]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_raddr_0[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0 [4])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_raddr_0<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_raddr_0[4]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_raddr_0[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18206.INIT = 16'hF0AA;
    X_LUT4 C18206(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2624 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/conf_latency_tim_out [6]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N42 )
    );
    defparam C18205.INIT = 16'hEE44;
    X_LUT4 C18205(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2625 ),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_latency_tim_out [7]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N48 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer_reg<6> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N42 ),
      .CLK (CLK_BUFGPed),
      .CE (N12351),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [6])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer_reg<7> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C2705/N48 ),
      .CLK (CLK_BUFGPed),
      .CE (N12351),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [7])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer[7]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18074.INIT = 16'hFAEA;
    X_LUT4 C18074(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/write_req_int ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/rdy_out358 )
    );
    defparam C19402.INIT = 16'h0004;
    X_LUT4 C19402(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/err_recovery ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .O (\bridge/wishbone_slave_unit/pcim_if_rdy_out/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_rdy_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_rdy_out/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_rdy_out/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_rdy_out/FROM ),
      .O (syn60010)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/rdy_out_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/rdy_out358 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/pcim_if_rdy_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_rdy_out )
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_rdy_out/FFY/ASYNC_FF_GSR_OR_6 (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_rdy_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_rdy_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17708.INIT = 16'h6666;
    X_LUT4 C17708(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [1]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [0]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [0])
    );
    defparam C17704.INIT = 16'h6666;
    X_LUT4 C17704(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [1]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [1])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [0])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<1>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [1])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<1>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17913.INIT = 16'h0011;
    X_LUT4 C17913(
      .ADR0 (\bridge/pci_target_unit/pcit_if_norm_access_to_config_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/req_comp_pending ),
      .O (\bridge/pci_target_unit/pci_target_sm/read_request )
    );
    defparam C17916.INIT = 16'hF5F0;
    X_LUT4 C17916(
      .ADR0 (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pcit_if_norm_access_to_config_out ),
      .ADR3 (syn19927),
      .O (\bridge/pci_target_unit/pci_target_sm/write_progress )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/wr_progress/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/wr_progress/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/rd_request_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/read_request ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/wr_progress/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/rd_request )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/wr_progress/FFY/ASYNC_FF_GSR_OR_7 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/wr_progress/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/wr_progress/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/wr_progress_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/write_progress ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/wr_progress/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/wr_progress )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/wr_progress/FFX/ASYNC_FF_GSR_OR_8 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/wr_progress/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/wr_progress/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17707.INIT = 16'h6666;
    X_LUT4 C17707(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [3]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [2])
    );
    defparam C17705.INIT = 16'h33CC;
    X_LUT4 C17705(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [3]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [4]),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [3])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [2])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<3>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [3])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<3>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17709.INIT = 16'h5A5A;
    X_LUT4 C17709(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [5]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [4]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [4])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_rgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [4])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<5>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next_reg<5> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [5])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<5>/FFX/SETOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFX/SET )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFX/SET ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next[5]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17618.INIT = 16'h5AAA;
    X_LUT4 C17618(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N361 )
    );
    defparam C17644.INIT = 16'h6CCC;
    X_LUT4 C17644(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N362 )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N361 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N362 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17660.INIT = 16'h3CCC;
    X_LUT4 C17660(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [0]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [1]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N345 )
    );
    defparam C17682.INIT = 16'h78F0;
    X_LUT4 C17682(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [0]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N346 )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N345 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N346 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17700.INIT = 16'h6A6A;
    X_LUT4 C17700(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [2])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [0])
      ,
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [1])
      ,
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N272 )
    );
    defparam C17714.INIT = 16'h6CCC;
    X_LUT4 C17714(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [0])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [3])
      ,
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [2])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [1])
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N273 )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N272 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [2])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<3>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N273 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [3])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<3>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17732.INIT = 16'h3CCC;
    X_LUT4 C17732(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [2])
      ,
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [1])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [0])
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N327 )
    );
    defparam C17754.INIT = 16'h7F80;
    X_LUT4 C17754(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [0])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [1])
      ,
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [2])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [3])
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N328 )
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one<3>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N327 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N328 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19477.INIT = 16'h2200;
    X_LUT4 C19477(
      .ADR0 (syn18858),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .ADR2 (VCC),
      .ADR3 (syn18863),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/GROM )
    );
    defparam C19474.INIT = 16'h0080;
    X_LUT4 C19474(
      .ADR0 (\bridge/in_reg_frame_out ),
      .ADR1 (\bridge/in_reg_irdy_out ),
      .ADR2 (N12359),
      .ADR3 (N_GNT),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<1>/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/GROM ),
      .O (N12359)
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/FROM ),
      .O (syn18937)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state_reg<1> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17620.INIT = 16'h3CF0;
    X_LUT4 C17620(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/C355/C3/C1 ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N363 )
    );
    defparam C17645.INIT = 16'h8080;
    X_LUT4 C17645(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [2]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<4>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/C355/C3/C1 )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N363 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<4>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[4]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17662.INIT = 16'h3CF0;
    X_LUT4 C17662(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/C333/C3/C1 ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N347 )
    );
    defparam C17683.INIT = 16'hC000;
    X_LUT4 C17683(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [0]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [1]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[4]/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one<4>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[4]/FROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/C333/C3/C1 )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N347 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[4]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[4]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17702.INIT = 16'h3C3C;
    X_LUT4 C17702(
      .ADR0 (VCC),
      .ADR1 (syn23402),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [4])
      ,
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N274 )
    );
    defparam C19443.INIT = 16'hF000;
    X_LUT4 C19443(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [4])
      ,
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FROM )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<4>/XUSED (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FROM ),
      .O (syn18958)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N274 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [4])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<4>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[4]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17734.INIT = 16'h66AA;
    X_LUT4 C17734(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [4])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [3])
      ,
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/C311/C3/C1 ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N329 )
    );
    defparam C17755.INIT = 16'h8080;
    X_LUT4 C17755(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [2])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [0])
      ,
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [1])
      ,
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FROM )
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<4>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/SRNOT )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<4>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FROM )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/C311/C3/C1 )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N329 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<4>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[4]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19469.INIT = 16'hF3F0;
    X_LUT4 C19469(
      .ADR0 (VCC),
      .ADR1 (\bridge/out_bckp_frame_out ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/GROM )
    );
    defparam C19484.INIT = 16'h0010;
    X_LUT4 C19484(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [0]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [2]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<2>/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C4/N9 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<2>/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state_reg<2> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[2]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17710.INIT = 16'h3CF0;
    X_LUT4 C17710(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [4])
      ,
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [5])
      ,
      .ADR3 (syn23402),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N275 )
    );
    defparam C17711.INIT = 16'h8000;
    X_LUT4 C17711(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [2])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [1])
      ,
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [0])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [3])
      ,
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FROM )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<5>/XUSED (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FROM ),
      .O (syn23402)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one_reg<5> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N275 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [5])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<5>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[5]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17934.INIT = 16'h5A5A;
    X_LUT4 C17934(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [1]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [0]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[0]/GROM )
    );
    X_INV \bridge/pci_target_unit/fifos/inGreyCount<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[0]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/inGreyCount<0>/YUSED (
      .I (\bridge/pci_target_unit/fifos/inGreyCount[0]/GROM ),
      .O (\bridge/pci_target_unit/fifos/inNextGreyCount [0])
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_inTransactionCount_reg<1> (
      .I (\bridge/pci_target_unit/fifos/inGreyCount[0]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/in_count_en ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/inGreyCount[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [1])
    );
    X_OR2 \bridge/pci_target_unit/fifos/inGreyCount<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/inGreyCount[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[0]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/inGreyCount_reg<0> (
      .I (\bridge/pci_target_unit/fifos/inNextGreyCount [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/in_count_en ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/inGreyCount[0]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/inGreyCount [0])
    );
    X_OR2 \bridge/pci_target_unit/fifos/inGreyCount<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/inGreyCount[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[0]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18215.INIT = 16'hC0C0;
    X_LUT4 C18215(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/out_bckp_frame_out ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C3/N5 )
    );
    defparam C19466.INIT = 16'hCC80;
    X_LUT4 C19466(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/out_bckp_frame_out ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<3>/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/FROM ),
      .O (syn18899)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state_reg<3> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C3/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[3]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17921.INIT = 16'h3FC0;
    X_LUT4 C17921(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [0]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [2]),
      .O (\bridge/pci_target_unit/fifos/N1961 )
    );
    defparam C17920.INIT = 16'h6CCC;
    X_LUT4 C17920(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [0]),
      .O (\bridge/pci_target_unit/fifos/N1962 )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_inTransactionCount<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_inTransactionCount_reg<2> (
      .I (\bridge/pci_target_unit/fifos/N1961 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/in_count_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_inTransactionCount<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_inTransactionCount_reg<3> (
      .I (\bridge/pci_target_unit/fifos/N1962 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/in_count_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_inTransactionCount<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17937.INIT = 16'hF050;
    X_LUT4 C17937(
      .ADR0 (\bridge/pci_target_unit/pcit_if_norm_access_to_config_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/conf_pci_img_ctrl1_out [0]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/decoder1/S_37/cell0 ),
      .O (\bridge/pci_target_unit/pci_target_if/C19/N5 )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C121 .INIT = 16'hAAA8;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C121 (
      .ADR0 (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_norm_access_to_config_out ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/config_access ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/decoder1/S_37/cell0 ),
      .O (\bridge/pciu_conf_offset_out[8]/FROM )
    );
    X_INV \bridge/pciu_conf_offset_out<8>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_conf_offset_out[8]/SRNOT )
    );
    X_BUF \bridge/pciu_conf_offset_out<8>/XUSED (
      .I (\bridge/pciu_conf_offset_out[8]/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn51 )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_prf_en_reg (
      .I (\bridge/pci_target_unit/pci_target_if/C19/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pciu_conf_offset_out[8]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/norm_prf_en )
    );
    X_OR2 \bridge/pciu_conf_offset_out<8>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_conf_offset_out[8]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_conf_offset_out[8]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<8> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pciu_conf_offset_out[8]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_conf_offset_out [8])
    );
    X_OR2 \bridge/pciu_conf_offset_out<8>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_conf_offset_out[8]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_conf_offset_out[8]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19356.INIT = 16'hC000;
    X_LUT4 C19356(
      .ADR0 (VCC),
      .ADR1 (N12360),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [10]),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/GROM )
    );
    defparam C19357.INIT = 16'hA000;
    X_LUT4 C19357(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [11]),
      .ADR1 (VCC),
      .ADR2 (N12360),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<11>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [10])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<11>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [11])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<10> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [10])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<11> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [11])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19417.INIT = 16'hC000;
    X_LUT4 C19417(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [20]),
      .ADR2 (syn24500),
      .ADR3 (N12360),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/GROM )
    );
    defparam C19418.INIT = 16'hA000;
    X_LUT4 C19418(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [21]),
      .ADR1 (VCC),
      .ADR2 (N12360),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<21>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [20])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<21>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [21])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<20> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [20])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<21> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [21])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[21]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19358.INIT = 16'hC000;
    X_LUT4 C19358(
      .ADR0 (VCC),
      .ADR1 (syn24500),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [12]),
      .ADR3 (N12360),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/GROM )
    );
    defparam C19359.INIT = 16'h8080;
    X_LUT4 C19359(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [13]),
      .ADR1 (N12360),
      .ADR2 (syn24500),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<13>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [12])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<13>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [13])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<12> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [12])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<13> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [13])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19427.INIT = 16'h8080;
    X_LUT4 C19427(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [30]),
      .ADR1 (N12360),
      .ADR2 (syn24500),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/GROM )
    );
    defparam C19428.INIT = 16'h8800;
    X_LUT4 C19428(
      .ADR0 (N12360),
      .ADR1 (syn24500),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [31]),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<31>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [30])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<31>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [31])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<30> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [30])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<31> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [31])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[31]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19419.INIT = 16'h8800;
    X_LUT4 C19419(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [22]),
      .ADR1 (N12360),
      .ADR2 (VCC),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/GROM )
    );
    defparam C19420.INIT = 16'h8800;
    X_LUT4 C19420(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [23]),
      .ADR1 (N12360),
      .ADR2 (VCC),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<23>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [22])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<23>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [23])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<22> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [22])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<23> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [23])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[23]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19360.INIT = 16'h8800;
    X_LUT4 C19360(
      .ADR0 (N12360),
      .ADR1 (syn24500),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [14]),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/GROM )
    );
    defparam C19361.INIT = 16'h8800;
    X_LUT4 C19361(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [15]),
      .ADR2 (VCC),
      .ADR3 (N12360),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<15>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [14])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<15>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [15])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<14> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [14])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<15> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [15])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19421.INIT = 16'hA000;
    X_LUT4 C19421(
      .ADR0 (syn24500),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [24]),
      .ADR3 (N12360),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/GROM )
    );
    defparam C19422.INIT = 16'hC000;
    X_LUT4 C19422(
      .ADR0 (VCC),
      .ADR1 (N12360),
      .ADR2 (syn24500),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [25]),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<25>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [24])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<25>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [25])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<24> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [24])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<25> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [25])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[25]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19413.INIT = 16'hA000;
    X_LUT4 C19413(
      .ADR0 (N12360),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [16]),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/GROM )
    );
    defparam C19414.INIT = 16'h8800;
    X_LUT4 C19414(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [17]),
      .ADR1 (syn24500),
      .ADR2 (VCC),
      .ADR3 (N12360),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<17>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [16])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<17>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [17])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<16> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [16])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<17> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [17])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17665.INIT = 16'hEECC;
    X_LUT4 C17665(
      .ADR0 (syn182579),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0 ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_almost_full_in )
    );
    defparam C17670.INIT = 16'hFCCC;
    X_LUT4 C17670(
      .ADR0 (VCC),
      .ADR1 (syn23568),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0 ),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_full )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/almost_full_reg (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_almost_full_in ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos_pcir_full_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/almost_full )
    );
    X_BUF \bridge/pci_target_unit/fifos_pcir_full_out/FFY/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos_pcir_full_out/FFY/RST )
    );
    X_OR2 \bridge/pci_target_unit/fifos_pcir_full_out/FFY/ASYNC_FF_GSR_OR_9 (
      .I0 (\bridge/pci_target_unit/fifos_pcir_full_out/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos_pcir_full_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/full_reg (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_full ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos_pcir_full_out/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos_pcir_full_out )
    );
    X_BUF \bridge/pci_target_unit/fifos_pcir_full_out/FFX/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos_pcir_full_out/FFX/RST )
    );
    X_OR2 \bridge/pci_target_unit/fifos_pcir_full_out/FFX/ASYNC_FF_GSR_OR_10 (
      .I0 (\bridge/pci_target_unit/fifos_pcir_full_out/FFX/RST ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos_pcir_full_out/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19423.INIT = 16'hA000;
    X_LUT4 C19423(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [26]),
      .ADR1 (VCC),
      .ADR2 (N12360),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/GROM )
    );
    defparam C19424.INIT = 16'h8080;
    X_LUT4 C19424(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [27]),
      .ADR1 (syn24500),
      .ADR2 (N12360),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<27>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [26])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<27>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [27])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<26> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [26])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<27> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [27])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[27]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19415.INIT = 16'h8800;
    X_LUT4 C19415(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [18]),
      .ADR2 (VCC),
      .ADR3 (N12360),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/GROM )
    );
    defparam C19416.INIT = 16'hC000;
    X_LUT4 C19416(
      .ADR0 (VCC),
      .ADR1 (syn24500),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [19]),
      .ADR3 (N12360),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<19>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [18])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<19>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [19])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<18> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [18])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<19> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [19])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17751.INIT = 16'h3C3C;
    X_LUT4 C17751(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [1]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [0]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next [0])
    );
    defparam C17736.INIT = 16'h0FF0;
    X_LUT4 C17736(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [1]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [2]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next [1])
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18066.INIT = 16'h5050;
    X_LUT4 C18066(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [0]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N192 )
    );
    defparam C18065.INIT = 16'h2222;
    X_LUT4 C18065(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [1]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N186 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<1>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<0> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N192 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<1> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N186 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17770.INIT = 16'h8888;
    X_LUT4 C17770(
      .ADR0 (\bridge/pci_target_unit/del_sync/N1245 ),
      .ADR1 (syn23138),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N55 )
    );
    defparam C17769.INIT = 16'h8888;
    X_LUT4 C17769(
      .ADR0 (syn23138),
      .ADR1 (\bridge/pci_target_unit/del_sync/N1246 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N60 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[11]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<10> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N55 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [10])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<11> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N60 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [11])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19425.INIT = 16'hC000;
    X_LUT4 C19425(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [28]),
      .ADR2 (N12360),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/GROM )
    );
    defparam C19426.INIT = 16'hC000;
    X_LUT4 C19426(
      .ADR0 (VCC),
      .ADR1 (N12360),
      .ADR2 (syn24500),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [29]),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_addr_out<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<29>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [28])
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_addr_out<29>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_data_out [29])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<28> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [28])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/addr_out_reg<29> (
      .I (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_addr_out [29])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_addr_out<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_addr_out[29]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18100.INIT = 16'h8888;
    X_LUT4 C18100(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/N150 ),
      .ADR1 (syn22149),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N55 )
    );
    defparam C18099.INIT = 16'hCC00;
    X_LUT4 C18099(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/N151 ),
      .ADR2 (VCC),
      .ADR3 (syn22149),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N60 )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<10> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N55 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [10])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<11> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N60 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/FFX/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [11])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17750.INIT = 16'h5A5A;
    X_LUT4 C17750(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [3]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [2]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next [2])
    );
    defparam C17741.INIT = 16'h5A5A;
    X_LUT4 C17741(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [3]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [4]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next [3])
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_rgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18064.INIT = 16'h4444;
    X_LUT4 C18064(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N180 )
    );
    defparam C18063.INIT = 16'h0A0A;
    X_LUT4 C18063(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [3]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N174 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<3>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<2> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N180 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<3> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N174 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17768.INIT = 16'h8888;
    X_LUT4 C17768(
      .ADR0 (\bridge/pci_target_unit/del_sync/N1247 ),
      .ADR1 (syn23138),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N65 )
    );
    defparam C17767.INIT = 16'h8888;
    X_LUT4 C17767(
      .ADR0 (syn23138),
      .ADR1 (\bridge/pci_target_unit/del_sync/N1248 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N70 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[13]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<12> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N65 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [12])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<13> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N70 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [13])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[13]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17938.INIT = 16'h8800;
    X_LUT4 C17938(
      .ADR0 (syn182016),
      .ADR1 (syn182017),
      .ADR2 (VCC),
      .ADR3 (syn182021),
      .O (\bridge/pci_target_unit/pci_target_sm/same_read_reg/GROM )
    );
    defparam C17939.INIT = 16'h8000;
    X_LUT4 C17939(
      .ADR0 (syn182005),
      .ADR1 (syn182015),
      .ADR2 (syn182004),
      .ADR3 (syn182018),
      .O (\bridge/pci_target_unit/pci_target_sm/same_read_reg/FROM )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/same_read_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/same_read_reg/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/same_read_reg/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/same_read_reg/GROM ),
      .O (N12467)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/same_read_reg/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/same_read_reg/FROM ),
      .O (syn182021)
    );
    X_FF \bridge/pci_target_unit/pci_target_if/same_read_reg_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/same_read_reg/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/same_read_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/same_read_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/same_read_reg/FFY/ASYNC_FF_GSR_OR_11 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/same_read_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/same_read_reg/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/same_read_reg_reg (
      .I (N12467),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/same_read_reg/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/same_read_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/same_read_reg/FFX/ASYNC_FF_GSR_OR_12 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/same_read_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/same_read_reg/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18098.INIT = 16'h8888;
    X_LUT4 C18098(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/N152 ),
      .ADR1 (syn22149),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N65 )
    );
    defparam C18097.INIT = 16'hC0C0;
    X_LUT4 C18097(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/N153 ),
      .ADR2 (syn22149),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N70 )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<12> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N65 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [12])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<13> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N70 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/FFX/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [13])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[13]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18062.INIT = 16'h0A0A;
    X_LUT4 C18062(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [4]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N168 )
    );
    defparam C18061.INIT = 16'h0A0A;
    X_LUT4 C18061(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [5]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N162 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<5>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<4> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N168 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<5> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N162 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [5])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[5]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17766.INIT = 16'hA0A0;
    X_LUT4 C17766(
      .ADR0 (\bridge/pci_target_unit/del_sync/N1249 ),
      .ADR1 (VCC),
      .ADR2 (syn23138),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N75 )
    );
    defparam C17765.INIT = 16'hC0C0;
    X_LUT4 C17765(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/N1250 ),
      .ADR2 (syn23138),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N80 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[15]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<14> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N75 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [14])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<15> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N80 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [15])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[15]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18096.INIT = 16'hAA00;
    X_LUT4 C18096(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/N154 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn22149),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N75 )
    );
    defparam C18095.INIT = 16'hCC00;
    X_LUT4 C18095(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/N155 ),
      .ADR2 (VCC),
      .ADR3 (syn22149),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N80 )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<14> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N75 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [14])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<15> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N80 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/FFX/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [15])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[15]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18961.INIT = 16'h5454;
    X_LUT4 C18961(
      .ADR0 (N12119),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbs_if/N40 )
    );
    defparam C18962.INIT = 16'h0200;
    X_LUT4 C18962(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR1 (ADR_O[2]),
      .ADR2 (ADR_O[10]),
      .ADR3 (N12119),
      .O (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FROM ),
      .O (N12118)
    );
    X_FF \CRT/ssvga_wbs_if/wbs_err_o_reg (
      .I (\CRT/ssvga_wbs_if/N40 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FFY/ASYNC_FF_GSR_OR ),
      .O (ERR_I)
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FFY/ASYNC_FF_GSR_OR_13 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF
     \bridge/wishbone_slave_unit/del_sync/rty_exp_sync/sync_data_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FFX/ASYNC_FF_GSR_OR_14 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18060.INIT = 16'h00AA;
    X_LUT4 C18060(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [6]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N156 )
    );
    defparam C18059.INIT = 16'h00CC;
    X_LUT4 C18059(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [7]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N150 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<7>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<6> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N156 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [6])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<7> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N150 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [7])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[7]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17764.INIT = 16'hF000;
    X_LUT4 C17764(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn23138),
      .ADR3 (\bridge/pci_target_unit/del_sync/N1251 ),
      .O (\bridge/pci_target_unit/del_sync/C1265/N85 )
    );
    defparam C17779.INIT = 16'hCC00;
    X_LUT4 C17779(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/N1236 ),
      .ADR2 (VCC),
      .ADR3 (syn23138),
      .O (\bridge/pci_target_unit/del_sync/C1265/N10 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<16> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N85 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [16])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<1> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N10 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [1])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18094.INIT = 16'h8888;
    X_LUT4 C18094(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/N156 ),
      .ADR1 (syn22149),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N85 )
    );
    defparam C18109.INIT = 16'hCC00;
    X_LUT4 C18109(
      .ADR0 (VCC),
      .ADR1 (syn22149),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/N141 ),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N10 )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<16> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N85 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [16])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<1> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N10 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18058.INIT = 16'h00AA;
    X_LUT4 C18058(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [8]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N144 )
    );
    defparam C18057.INIT = 16'h00CC;
    X_LUT4 C18057(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [9]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N138 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<9>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<8> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N144 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [8])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<9> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N138 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [9])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[9]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17890.INIT = 16'hFF88;
    X_LUT4 C17890(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [0]),
      .ADR1 (syn16925),
      .ADR2 (VCC),
      .ADR3 (syn182122),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N6 )
    );
    defparam C17891.INIT = 16'hD5C0;
    X_LUT4 C17891(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [0]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N2983 ),
      .O (\bridge/pciu_err_addr_out[0]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[0]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<0>/XUSED (
      .I (\bridge/pciu_err_addr_out[0]/FROM ),
      .O (syn182122)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<0> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[0] )
    );
    X_OR2 \bridge/pciu_err_addr_out<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18140.INIT = 16'hBBBB;
    X_LUT4 C18140(
      .ADR0 (\bridge/conf_wb_err_pending_out ),
      .ADR1 (\bridge/conf_pci_master_enable_out ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/wbs_sm_lock_in )
    );
    defparam C19511.INIT = 16'hECA0;
    X_LUT4 C19511(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [2]),
      .ADR1 (syn24559),
      .ADR2 (syn17745),
      .ADR3 (\bridge/conf_pci_master_enable_out ),
      .O (\bridge/in_reg_idsel_out/FROM )
    );
    X_INV \bridge/in_reg_idsel_out/SRMUX (
      .I (N_RST),
      .O (\bridge/in_reg_idsel_out/SRNOT )
    );
    X_BUF \bridge/in_reg_idsel_out/XUSED (
      .I (\bridge/in_reg_idsel_out/FROM ),
      .O (syn178469)
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/lock_reg (
      .I (\bridge/wishbone_slave_unit/wbs_sm_lock_in ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/in_reg_idsel_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/lock )
    );
    X_OR2 \bridge/in_reg_idsel_out/FFY/ASYNC_FF_GSR_OR_15 (
      .I0 (\bridge/in_reg_idsel_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/in_reg_idsel_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/input_register/pci_idsel_reg_out_reg (
      .I (N_IDSEL),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/in_reg_idsel_out/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/in_reg_idsel_out )
    );
    X_OR2 \bridge/in_reg_idsel_out/FFX/ASYNC_FF_GSR_OR_16 (
      .I0 (\bridge/in_reg_idsel_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/in_reg_idsel_out/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17887.INIT = 16'hFF88;
    X_LUT4 C17887(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [1]),
      .ADR1 (syn16925),
      .ADR2 (VCC),
      .ADR3 (syn182129),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N12 )
    );
    defparam C17888.INIT = 16'hCE0A;
    X_LUT4 C17888(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N2984 ),
      .ADR1 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [1]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR3 (syn16933),
      .O (\bridge/pciu_err_addr_out[1]/FROM )
    );
    X_INV \bridge/pciu_err_addr_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_addr_out[1]/SRNOT )
    );
    X_BUF \bridge/pciu_err_addr_out<1>/XUSED (
      .I (\bridge/pciu_err_addr_out[1]/FROM ),
      .O (syn182129)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<1> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\bridge/pciu_err_addr_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_addr_out[1] )
    );
    X_OR2 \bridge/pciu_err_addr_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_addr_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_addr_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17885.INIT = 16'hFFC0;
    X_LUT4 C17885(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [2]),
      .ADR2 (syn16925),
      .ADR3 (syn182134),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N18 )
    );
    defparam C17886.INIT = 16'h88F8;
    X_LUT4 C17886(
      .ADR0 (syn16933),
      .ADR1 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [2]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/N2985 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\ADR_O[2]/FROM )
    );
    X_INV \ADR_O<2>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[2]/SRNOT )
    );
    X_BUF \ADR_O<2>/XUSED (
      .I (\ADR_O[2]/FROM ),
      .O (syn182134)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<2> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[2]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[2])
    );
    X_OR2 \ADR_O<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[2]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[2]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C20039.INIT = 16'hF0CC;
    X_LUT4 C20039(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_be_out [2]),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_cbe_out [2]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .O (\bridge/configuration/pci_err_cs_bit31_24[30]/GROM )
    );
    defparam C20040.INIT = 16'h000A;
    X_LUT4 C20040(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/c_state [0]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/c_state [1]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/c_state [2]),
      .O (\bridge/configuration/pci_err_cs_bit31_24[30]/FROM )
    );
    X_INV \bridge/configuration/pci_err_cs_bit31_24<30>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_cs_bit31_24[30]/SRNOT )
    );
    X_BUF \bridge/configuration/pci_err_cs_bit31_24<30>/YUSED (
      .I (\bridge/configuration/pci_err_cs_bit31_24[30]/GROM ),
      .O (N12519)
    );
    X_BUF \bridge/configuration/pci_err_cs_bit31_24<30>/XUSED (
      .I (\bridge/configuration/pci_err_cs_bit31_24[30]/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C981 )
    );
    X_FF \bridge/configuration/pci_err_cs_bit31_24_reg<30> (
      .I (\bridge/configuration/pci_err_cs_bit31_24[30]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_cs_bit31_24[30]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_cs_bit31_24 [30])
    );
    X_OR2 \bridge/configuration/pci_err_cs_bit31_24<30>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_cs_bit31_24[30]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_cs_bit31_24[30]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17883.INIT = 16'hFF88;
    X_LUT4 C17883(
      .ADR0 (syn16925),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [3]),
      .ADR2 (VCC),
      .ADR3 (syn182139),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N24 )
    );
    defparam C17884.INIT = 16'hB3A0;
    X_LUT4 C17884(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [3]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR2 (syn16933),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N2986 ),
      .O (\ADR_O[3]/FROM )
    );
    X_INV \ADR_O<3>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[3]/SRNOT )
    );
    X_BUF \ADR_O<3>/XUSED (
      .I (\ADR_O[3]/FROM ),
      .O (syn182139)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<3> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N24 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[3])
    );
    X_OR2 \ADR_O<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[3]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[3]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18814.INIT = 16'hE2E2;
    X_LUT4 C18814(
      .ADR0 (\bridge/pci_target_unit/del_sync_be_out [3]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_cbe_out [3]),
      .ADR3 (VCC),
      .O (N12518)
    );
    defparam C18960.INIT = 16'h2000;
    X_LUT4 C18960(
      .ADR0 (N12119),
      .ADR1 (ADR_O[10]),
      .ADR2 (ADR_O[2]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .O (\bridge/configuration/pci_err_cs_bit31_24[31]/FROM )
    );
    X_INV \bridge/configuration/pci_err_cs_bit31_24<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_cs_bit31_24[31]/SRNOT )
    );
    X_BUF \bridge/configuration/pci_err_cs_bit31_24<31>/XUSED (
      .I (\bridge/configuration/pci_err_cs_bit31_24[31]/FROM ),
      .O (N12120)
    );
    X_FF \bridge/configuration/pci_err_cs_bit31_24_reg<31> (
      .I (N12518),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_cs_bit31_24[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_cs_bit31_24 [31])
    );
    X_OR2 \bridge/configuration/pci_err_cs_bit31_24<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_cs_bit31_24[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_cs_bit31_24[31]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17881.INIT = 16'hFFA0;
    X_LUT4 C17881(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [4]),
      .ADR1 (VCC),
      .ADR2 (syn16925),
      .ADR3 (syn182144),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N30 )
    );
    defparam C17882.INIT = 16'hAE0C;
    X_LUT4 C17882(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [4]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N2987 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR3 (syn16933),
      .O (\ADR_O[4]/FROM )
    );
    X_INV \ADR_O<4>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[4]/SRNOT )
    );
    X_BUF \ADR_O<4>/XUSED (
      .I (\ADR_O[4]/FROM ),
      .O (syn182144)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<4> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[4])
    );
    X_OR2 \ADR_O<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[4]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17879.INIT = 16'hFF88;
    X_LUT4 C17879(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [5]),
      .ADR1 (syn16925),
      .ADR2 (VCC),
      .ADR3 (syn182149),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N36 )
    );
    defparam C17880.INIT = 16'hD5C0;
    X_LUT4 C17880(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [5]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N2988 ),
      .O (\ADR_O[5]/FROM )
    );
    X_INV \ADR_O<5>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[5]/SRNOT )
    );
    X_BUF \ADR_O<5>/XUSED (
      .I (\ADR_O[5]/FROM ),
      .O (syn182149)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<5> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[5])
    );
    X_OR2 \ADR_O<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[5]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[5]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17877.INIT = 16'hFF88;
    X_LUT4 C17877(
      .ADR0 (syn16925),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [6]),
      .ADR2 (VCC),
      .ADR3 (syn182154),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N42 )
    );
    defparam C17878.INIT = 16'hD5C0;
    X_LUT4 C17878(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [6]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N2989 ),
      .O (\ADR_O[6]/FROM )
    );
    X_INV \ADR_O<6>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[6]/SRNOT )
    );
    X_BUF \ADR_O<6>/XUSED (
      .I (\ADR_O[6]/FROM ),
      .O (syn182154)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<6> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N42 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[6]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[6])
    );
    X_OR2 \ADR_O<6>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[6]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[6]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17875.INIT = 16'hFFC0;
    X_LUT4 C17875(
      .ADR0 (VCC),
      .ADR1 (syn16925),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [7]),
      .ADR3 (syn182159),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N48 )
    );
    defparam C17876.INIT = 16'hC0EA;
    X_LUT4 C17876(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N2990 ),
      .ADR1 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [7]),
      .ADR2 (syn16933),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\ADR_O[7]/FROM )
    );
    X_INV \ADR_O<7>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[7]/SRNOT )
    );
    X_BUF \ADR_O<7>/XUSED (
      .I (\ADR_O[7]/FROM ),
      .O (syn182159)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<7> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N48 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[7])
    );
    X_OR2 \ADR_O<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[7]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[7]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17873.INIT = 16'hFF88;
    X_LUT4 C17873(
      .ADR0 (syn16925),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [8]),
      .ADR2 (VCC),
      .ADR3 (syn182164),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N54 )
    );
    defparam C17874.INIT = 16'hB3A0;
    X_LUT4 C17874(
      .ADR0 (syn16933),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [8]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N2991 ),
      .O (\ADR_O[8]/FROM )
    );
    X_INV \ADR_O<8>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[8]/SRNOT )
    );
    X_BUF \ADR_O<8>/XUSED (
      .I (\ADR_O[8]/FROM ),
      .O (syn182164)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<8> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N54 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[8]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[8])
    );
    X_OR2 \ADR_O<8>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[8]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[8]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C20038.INIT = 16'hFA50;
    X_LUT4 C20038(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync_be_out [0]),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_cbe_out [0]),
      .O (\bridge/configuration/pci_err_cs_bit31_24[29]/GROM )
    );
    defparam C20037.INIT = 16'hEE44;
    X_LUT4 C20037(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR1 (\bridge/pci_target_unit/del_sync_be_out [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_cbe_out [1]),
      .O (\bridge/configuration/pci_err_cs_bit31_24[29]/FROM )
    );
    X_INV \bridge/configuration/pci_err_cs_bit31_24<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_cs_bit31_24[29]/SRNOT )
    );
    X_BUF \bridge/configuration/pci_err_cs_bit31_24<29>/YUSED (
      .I (\bridge/configuration/pci_err_cs_bit31_24[29]/GROM ),
      .O (N12521)
    );
    X_BUF \bridge/configuration/pci_err_cs_bit31_24<29>/XUSED (
      .I (\bridge/configuration/pci_err_cs_bit31_24[29]/FROM ),
      .O (N12520)
    );
    X_FF \bridge/configuration/pci_err_cs_bit31_24_reg<28> (
      .I (\bridge/configuration/pci_err_cs_bit31_24[29]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_cs_bit31_24[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_cs_bit31_24 [28])
    );
    X_OR2 \bridge/configuration/pci_err_cs_bit31_24<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_cs_bit31_24[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_cs_bit31_24[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_cs_bit31_24_reg<29> (
      .I (\bridge/configuration/pci_err_cs_bit31_24[29]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_cs_bit31_24[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_cs_bit31_24 [29])
    );
    X_OR2 \bridge/configuration/pci_err_cs_bit31_24<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_cs_bit31_24[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_cs_bit31_24[29]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17871.INIT = 16'hFF88;
    X_LUT4 C17871(
      .ADR0 (syn16925),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [9]),
      .ADR2 (VCC),
      .ADR3 (syn182169),
      .O (\bridge/pci_target_unit/wishbone_master/C3415/N60 )
    );
    defparam C17872.INIT = 16'hDC50;
    X_LUT4 C17872(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (syn16933),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/N2992 ),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_addr_data_out [9]),
      .O (\ADR_O[9]/FROM )
    );
    X_INV \ADR_O<9>/SRMUX (
      .I (N_RST),
      .O (\ADR_O[9]/SRNOT )
    );
    X_BUF \ADR_O<9>/XUSED (
      .I (\ADR_O[9]/FROM ),
      .O (syn182169)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/addr_cnt_out_reg<9> (
      .I (\bridge/pci_target_unit/wishbone_master/C3415/N60 ),
      .CLK (CLK_BUFGPed),
      .CE (N12478),
      .SET (GND),
      .RST (\ADR_O[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (ADR_O[9])
    );
    X_OR2 \ADR_O<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\ADR_O[9]/SRNOT ),
      .I1 (GSR),
      .O (\ADR_O[9]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17613.INIT = 16'h33CC;
    X_LUT4 C17613(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_waddr [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_waddr [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/GROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<0>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/GROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next [0])
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<0>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/waddr_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_waddr [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17611.INIT = 16'h5AAA;
    X_LUT4 C17611(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_waddr [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_waddr [0]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_waddr [1]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N322 )
    );
    defparam C17609.INIT = 16'h6AAA;
    X_LUT4 C17609(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_waddr [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_waddr [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_waddr [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_waddr [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N323 )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_waddr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[3]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_waddr<3>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[3]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/waddr_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N322 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_waddr[3]/CENOT ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_waddr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr [2])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_waddr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_waddr[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/waddr_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N323 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_waddr[3]/CENOT ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_waddr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr [3])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_waddr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_waddr[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17608.INIT = 16'h3CF0;
    X_LUT4 C17608(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_waddr [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_waddr [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/C354/C3/C1 ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N324 )
    );
    defparam C17610.INIT = 16'hC000;
    X_LUT4 C17610(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_waddr [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_waddr [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_waddr [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[4]/FROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_waddr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[4]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_waddr<4>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_waddr[4]/FROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/C354/C3/C1 )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_waddr<4>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[4]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/waddr_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N324 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_waddr[4]/CENOT ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_waddr[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr [4])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_waddr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_waddr[4]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17679.INIT = 16'h6666;
    X_LUT4 C17679(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [1]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next [0])
    );
    defparam C17664.INIT = 16'h6666;
    X_LUT4 C17664(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [1]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next [1])
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17678.INIT = 16'h0FF0;
    X_LUT4 C17678(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [3]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next [2])
    );
    defparam C17669.INIT = 16'h33CC;
    X_LUT4 C17669(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [4]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [3]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next [3])
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_rgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18266.INIT = 16'hFFA0;
    X_LUT4 C18266(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_bc_out [0]),
      .ADR3 (syn181290),
      .O (\bridge/out_bckp_cbe_out[0]/GROM )
    );
    defparam C18267.INIT = 16'hF888;
    X_LUT4 C18267(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_be_out [0]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_be_out [0]),
      .ADR3 (syn20493),
      .O (\bridge/out_bckp_cbe_out[0]/FROM )
    );
    X_INV \bridge/out_bckp_cbe_out<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_cbe_out[0]/SRNOT )
    );
    X_BUF \bridge/out_bckp_cbe_out<0>/YUSED (
      .I (\bridge/out_bckp_cbe_out[0]/GROM ),
      .O (\bridge/pci_mux_cbe_in [0])
    );
    X_BUF \bridge/out_bckp_cbe_out<0>/XUSED (
      .I (\bridge/out_bckp_cbe_out[0]/FROM ),
      .O (syn181290)
    );
    X_FF \bridge/output_backup/cbe_out_reg<0> (
      .I (\bridge/out_bckp_cbe_out[0]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_mas_load_in ),
      .SET (\bridge/out_bckp_cbe_out[0]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_cbe_out [0])
    );
    X_OR2 \bridge/out_bckp_cbe_out<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_cbe_out[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_cbe_out[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19143.INIT = 16'h0B0A;
    X_LUT4 C19143(
      .ADR0 (syn179287),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR2 (\bridge/in_reg_frame_out ),
      .ADR3 (syn19933),
      .O (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/GROM )
    );
    defparam C19146.INIT = 16'hFD5D;
    X_LUT4 C19146(
      .ADR0 (syn19407),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg [0]),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_control_out [0]),
      .O (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/FROM )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_disconect_wo_data_out )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/FROM ),
      .O (syn19933)
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/FFY/ASYNC_FF_GSR_OR_17 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C18261.INIT = 16'hFFA0;
    X_LUT4 C18261(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_bc_out [1]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR3 (syn181303),
      .O (\bridge/out_bckp_cbe_out[1]/GROM )
    );
    defparam C18262.INIT = 16'hEAC0;
    X_LUT4 C18262(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_be_out [1]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_be_out [1]),
      .O (\bridge/out_bckp_cbe_out[1]/FROM )
    );
    X_INV \bridge/out_bckp_cbe_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_cbe_out[1]/SRNOT )
    );
    X_BUF \bridge/out_bckp_cbe_out<1>/YUSED (
      .I (\bridge/out_bckp_cbe_out[1]/GROM ),
      .O (\bridge/pci_mux_cbe_in [1])
    );
    X_BUF \bridge/out_bckp_cbe_out<1>/XUSED (
      .I (\bridge/out_bckp_cbe_out[1]/FROM ),
      .O (syn181303)
    );
    X_FF \bridge/output_backup/cbe_out_reg<1> (
      .I (\bridge/out_bckp_cbe_out[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_mas_load_in ),
      .SET (\bridge/out_bckp_cbe_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_cbe_out [1])
    );
    X_OR2 \bridge/out_bckp_cbe_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_cbe_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_cbe_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C20020.INIT = 16'hFFCC;
    X_LUT4 C20020(
      .ADR0 (VCC),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/output_backup/mas_ad_en_out ),
      .O (\bridge/out_bckp_par_en_out/GROM )
    );
    X_INV \bridge/out_bckp_par_en_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_par_en_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_par_en_out/YUSED (
      .I (\bridge/out_bckp_par_en_out/GROM ),
      .O (\bridge/pci_mux_par_en_in )
    );
    X_FF \bridge/output_backup/par_en_out_reg (
      .I (\bridge/out_bckp_par_en_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/out_bckp_par_en_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_par_en_out )
    );
    X_OR2 \bridge/out_bckp_par_en_out/FFY/ASYNC_FF_GSR_OR_18 (
      .I0 (\bridge/out_bckp_par_en_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_par_en_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18256.INIT = 16'hFFA0;
    X_LUT4 C18256(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_bc_out [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR3 (syn181316),
      .O (\bridge/out_bckp_cbe_out[2]/GROM )
    );
    defparam C18257.INIT = 16'hECA0;
    X_LUT4 C18257(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_be_out [2]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_be_out [2]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .O (\bridge/out_bckp_cbe_out[2]/FROM )
    );
    X_INV \bridge/out_bckp_cbe_out<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_cbe_out[2]/SRNOT )
    );
    X_BUF \bridge/out_bckp_cbe_out<2>/YUSED (
      .I (\bridge/out_bckp_cbe_out[2]/GROM ),
      .O (\bridge/pci_mux_cbe_in [2])
    );
    X_BUF \bridge/out_bckp_cbe_out<2>/XUSED (
      .I (\bridge/out_bckp_cbe_out[2]/FROM ),
      .O (syn181316)
    );
    X_FF \bridge/output_backup/cbe_out_reg<2> (
      .I (\bridge/out_bckp_cbe_out[2]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_mas_load_in ),
      .SET (\bridge/out_bckp_cbe_out[2]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_cbe_out [2])
    );
    X_OR2 \bridge/out_bckp_cbe_out<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_cbe_out[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_cbe_out[2]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18251.INIT = 16'hFFC0;
    X_LUT4 C18251(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_bc_out [3]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR3 (syn181329),
      .O (\bridge/out_bckp_cbe_out[3]/GROM )
    );
    defparam C18252.INIT = 16'hF888;
    X_LUT4 C18252(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_be_out [3]),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_next_be_out [3]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .O (\bridge/out_bckp_cbe_out[3]/FROM )
    );
    X_INV \bridge/out_bckp_cbe_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_cbe_out[3]/SRNOT )
    );
    X_BUF \bridge/out_bckp_cbe_out<3>/YUSED (
      .I (\bridge/out_bckp_cbe_out[3]/GROM ),
      .O (\bridge/pci_mux_cbe_in [3])
    );
    X_BUF \bridge/out_bckp_cbe_out<3>/XUSED (
      .I (\bridge/out_bckp_cbe_out[3]/FROM ),
      .O (syn181329)
    );
    X_FF \bridge/output_backup/cbe_out_reg<3> (
      .I (\bridge/out_bckp_cbe_out[3]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_mas_load_in ),
      .SET (\bridge/out_bckp_cbe_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_cbe_out [3])
    );
    X_OR2 \bridge/out_bckp_cbe_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_cbe_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_cbe_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19259.INIT = 16'h0F0A;
    X_LUT4 C19259(
      .ADR0 (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out [1]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_full_out ),
      .ADR3 (syn17090),
      .O (\bridge/pci_target_unit/fifos/pcir_write_performed/GROM )
    );
    defparam C19260.INIT = 16'h0A00;
    X_LUT4 C19260(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .ADR1 (VCC),
      .ADR2 (ERR_I),
      .ADR3 (ACK_I),
      .O (\bridge/pci_target_unit/fifos/pcir_write_performed/FROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pcir_write_performed/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pcir_write_performed/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_write_performed/YUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_write_performed/GROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_wallow )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_write_performed/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_write_performed/FROM ),
      .O (syn17090)
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_write_performed_reg (
      .I (\bridge/pci_target_unit/fifos/pcir_write_performed/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_write_performed/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_write_performed )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_write_performed/FFY/ASYNC_FF_GSR_OR_19 (
      .I0 (\bridge/pci_target_unit/fifos/pcir_write_performed/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_write_performed/FFY/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_sm/frame_iob_en_feed/C40 .INIT = 16'hFF80;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_sm/frame_iob_en_feed/C40 (
      .ADR0 (N_STOP),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/frame_en_keep ),
      .ADR2 (N_TRDY),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/frame_en_slow ),
      .O (\bridge/out_bckp_frame_en_out/GROM )
    );
    defparam C19468.INIT = 16'hFFCE;
    X_LUT4 C19468(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (syn16939),
      .ADR2 (\bridge/out_bckp_frame_out ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .O (\bridge/out_bckp_frame_en_out/FROM )
    );
    X_INV \bridge/out_bckp_frame_en_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_frame_en_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_frame_en_out/YUSED (
      .I (\bridge/out_bckp_frame_en_out/GROM ),
      .O (\bridge/pci_mux_frame_en_in )
    );
    X_BUF \bridge/out_bckp_frame_en_out/XUSED (
      .I (\bridge/out_bckp_frame_en_out/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/frame_en_slow )
    );
    X_FF \bridge/output_backup/frame_en_out_reg (
      .I (\bridge/out_bckp_frame_en_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/out_bckp_frame_en_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_frame_en_out )
    );
    X_OR2 \bridge/out_bckp_frame_en_out/FFY/ASYNC_FF_GSR_OR_20 (
      .I0 (\bridge/out_bckp_frame_en_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_frame_en_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17803.INIT = 16'h00AA;
    X_LUT4 C17803(
      .ADR0 (syn17006),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [0]),
      .O (\bridge/pci_target_unit/wishbone_master/C103/N5 )
    );
    defparam C17801.INIT = 16'h2828;
    X_LUT4 C17801(
      .ADR0 (syn17006),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [0]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [1]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/C103/N10 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt_reg<0> (
      .I (\bridge/pci_target_unit/wishbone_master/C103/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/C104/N6 ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [0])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt_reg<1> (
      .I (\bridge/pci_target_unit/wishbone_master/C103/N10 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/C104/N6 ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [1])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19461.INIT = 16'hEEEE;
    X_LUT4 C19461(
      .ADR0 (syn18919),
      .ADR1 (syn178584),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_last_out )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_last_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_last_out/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/current_last_reg (
      .I (\bridge/wishbone_slave_unit/pcim_if_next_last_out ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/last_load ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/pcim_if_last_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_last_out )
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_last_out/FFY/ASYNC_FF_GSR_OR_21 (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_last_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_last_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18980.INIT = 16'hA0A0;
    X_LUT4 C18980(
      .ADR0 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr_plus1 [0]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C2/N50 )
    );
    defparam C18979.INIT = 16'hAA00;
    X_LUT4 C18979(
      .ADR0 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr_plus1 [1]),
      .O (\CRT/ssvga_fifo/C2/N45 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr[1]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<0> (
      .I (\CRT/ssvga_fifo/C2/N50 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [0])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<1> (
      .I (\CRT/ssvga_fifo/C2/N45 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [1])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19030.INIT = 16'hDD88;
    X_LUT4 C19030(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/pix_start_addr [2]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/N1717 ),
      .O (\CRT/ssvga_wbm_if/C1475/N6 )
    );
    defparam C19029.INIT = 16'hF5A0;
    X_LUT4 C19029(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [3]),
      .ADR3 (\CRT/ssvga_wbm_if/N1718 ),
      .O (\CRT/ssvga_wbm_if/C1475/N12 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<2> (
      .I (\CRT/ssvga_wbm_if/C1475/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2])
    );
    X_OR2 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<3> (
      .I (\CRT/ssvga_wbm_if/C1475/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3])
    );
    X_OR2 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18073.INIT = 16'h0300;
    X_LUT4 C18073(
      .ADR0 (VCC),
      .ADR1 (N_TRDY),
      .ADR2 (syn18863),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_last_out ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/last_transfered265 )
    );
    defparam C18222.INIT = 16'h0C0C;
    X_LUT4 C18222(
      .ADR0 (VCC),
      .ADR1 (syn21738),
      .ADR2 (syn18863),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout509 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/timeout/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/last_transfered_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/last_transfered265 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_control_out [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/timeout/FFY/ASYNC_FF_GSR_OR_22 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/timeout_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout509 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/timeout/FFX/ASYNC_FF_GSR_OR_23 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18075.INIT = 16'hCC00;
    X_LUT4 C18075(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [0]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C26/N6 )
    );
    defparam C18076.INIT = 16'hCCAA;
    X_LUT4 C18076(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_bc_out [1]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C26/N12 )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_bc_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/bc_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C26/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12594),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/pcim_if_bc_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out [0])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_bc_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_bc_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/bc_out_reg<1> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C26/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (N12594),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/pcim_if_bc_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out [1])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_bc_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_bc_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18978.INIT = 16'hAA00;
    X_LUT4 C18978(
      .ADR0 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr_plus1 [2]),
      .O (\CRT/ssvga_fifo/C2/N40 )
    );
    defparam C18977.INIT = 16'hA0A0;
    X_LUT4 C18977(
      .ADR0 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr_plus1 [3]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C2/N35 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr[3]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<2> (
      .I (\CRT/ssvga_fifo/C2/N40 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [2])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<3> (
      .I (\CRT/ssvga_fifo/C2/N35 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [3])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17797.INIT = 16'hA888;
    X_LUT4 C17797(
      .ADR0 (syn17006),
      .ADR1 (syn23094),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [3]),
      .ADR3 (syn23093),
      .O (\bridge/pci_target_unit/wishbone_master/C103/N20 )
    );
    defparam C17799.INIT = 16'h3FBF;
    X_LUT4 C17799(
      .ADR0 (syn17006),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [1]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [2]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [0]),
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/FROM )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<3>/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/FROM ),
      .O (syn23093)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt_reg<3> (
      .I (\bridge/pci_target_unit/wishbone_master/C103/N20 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/C104/N6 ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [3])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[3]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C19028.INIT = 16'hFA50;
    X_LUT4 C19028(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_wbm_if/N1719 ),
      .ADR3 (\CRT/pix_start_addr [4]),
      .O (\CRT/ssvga_wbm_if/C1475/N18 )
    );
    defparam C19027.INIT = 16'hACAC;
    X_LUT4 C19027(
      .ADR0 (\CRT/pix_start_addr [5]),
      .ADR1 (\CRT/ssvga_wbm_if/N1720 ),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1475/N24 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<4> (
      .I (\CRT/ssvga_wbm_if/C1475/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4])
    );
    X_OR2 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<5> (
      .I (\CRT/ssvga_wbm_if/C1475/N24 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5])
    );
    X_OR2 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18072.INIT = 16'hAAF0;
    X_LUT4 C18072(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_bc_out [2]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C26/N18 )
    );
    defparam C18080.INIT = 16'hEE22;
    X_LUT4 C18080(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_bc_out [3]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [3]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C26/N24 )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_bc_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/bc_out_reg<2> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C26/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (N12594),
      .SET (\bridge/wishbone_slave_unit/pcim_if_bc_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out [2])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_bc_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/bc_out_reg<3> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C26/N24 ),
      .CLK (CLK_BUFGPed),
      .CE (N12594),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/pcim_if_bc_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out [3])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_bc_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_bc_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18976.INIT = 16'hF000;
    X_LUT4 C18976(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr_plus1 [4]),
      .O (\CRT/ssvga_fifo/C2/N30 )
    );
    defparam C18975.INIT = 16'hF000;
    X_LUT4 C18975(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr_plus1 [5]),
      .ADR3 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .O (\CRT/ssvga_fifo/C2/N25 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr[5]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<4> (
      .I (\CRT/ssvga_fifo/C2/N30 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [4])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<5> (
      .I (\CRT/ssvga_fifo/C2/N25 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [5])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19026.INIT = 16'hDD88;
    X_LUT4 C19026(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/pix_start_addr [6]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/N1721 ),
      .O (\CRT/ssvga_wbm_if/C1475/N30 )
    );
    defparam C19025.INIT = 16'hFC30;
    X_LUT4 C19025(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR2 (\CRT/ssvga_wbm_if/N1722 ),
      .ADR3 (\CRT/pix_start_addr [7]),
      .O (\CRT/ssvga_wbm_if/C1475/N36 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<6> (
      .I (\CRT/ssvga_wbm_if/C1475/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6])
    );
    X_OR2 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<7> (
      .I (\CRT/ssvga_wbm_if/C1475/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7])
    );
    X_OR2 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18974.INIT = 16'hA0A0;
    X_LUT4 C18974(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr_plus1 [6]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C2/N20 )
    );
    defparam C18973.INIT = 16'hA0A0;
    X_LUT4 C18973(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr_plus1 [7]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C2/N15 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr[7]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<6> (
      .I (\CRT/ssvga_fifo/C2/N20 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [6])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<7> (
      .I (\CRT/ssvga_fifo/C2/N15 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [7])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19024.INIT = 16'hE2E2;
    X_LUT4 C19024(
      .ADR0 (\CRT/ssvga_wbm_if/N1723 ),
      .ADR1 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR2 (\CRT/pix_start_addr [8]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1475/N42 )
    );
    defparam C19023.INIT = 16'hEE22;
    X_LUT4 C19023(
      .ADR0 (\CRT/ssvga_wbm_if/N1724 ),
      .ADR1 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR2 (VCC),
      .ADR3 (\CRT/pix_start_addr [9]),
      .O (\CRT/ssvga_wbm_if/C1475/N48 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<8> (
      .I (\CRT/ssvga_wbm_if/C1475/N42 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [8])
    );
    X_OR2 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<9> (
      .I (\CRT/ssvga_wbm_if/C1475/N48 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [9])
    );
    X_OR2 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18972.INIT = 16'hCC00;
    X_LUT4 C18972(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [8]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .O (\CRT/ssvga_fifo/C2/N10 )
    );
    defparam C18971.INIT = 16'hC0C0;
    X_LUT4 C18971(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [9]),
      .ADR2 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C2/N5 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr<9>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr[9]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<8> (
      .I (\CRT/ssvga_fifo/C2/N10 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [8])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_reg<9> (
      .I (\CRT/ssvga_fifo/C2/N5 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr [9])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19963.INIT = 16'hCC00;
    X_LUT4 C19963(
      .ADR0 (VCC),
      .ADR1 (syn177380),
      .ADR2 (VCC),
      .ADR3 (syn177381),
      .O (\bridge/wishbone_slave_unit/amux_hit_out [1])
    );
    defparam C19964.INIT = 16'h8000;
    X_LUT4 C19964(
      .ADR0 (syn177391),
      .ADR1 (syn60044),
      .ADR2 (syn60045),
      .ADR3 (syn60043),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/wishbone_slave/img_hit<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/img_hit<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/FROM ),
      .O (syn177381)
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/img_hit_reg<0> (
      .I (\bridge/wishbone_slave_unit/amux_hit_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/img_hit [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/img_hit<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/img_hit[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17716.INIT = 16'hDD55;
    X_LUT4 C17716(
      .ADR0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect70 ),
      .ADR1 (syn182488),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/reg_empty )
    );
    defparam C19431.INIT = 16'hA0A0;
    X_LUT4 C19431(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [0])
      ,
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FROM ),
      .O (syn18984)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty_reg (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/reg_empty ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FFY/SETOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FFY/SET )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR_24 (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FFY/SET ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18998.INIT = 16'hBBBB;
    X_LUT4 C18998(
      .ADR0 (\CRT/ssvga_fifo/N738 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C751/N6 )
    );
    defparam C18981.INIT = 16'h8888;
    X_LUT4 C18981(
      .ADR0 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR1 (\CRT/ssvga_fifo/N739 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C751/N11 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr_plus1<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[1]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<0> (
      .I (\CRT/ssvga_fifo/C751/N6 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (\CRT/ssvga_fifo/rd_ptr_plus1[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [0])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<1> (
      .I (\CRT/ssvga_fifo/C751/N11 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [1])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18995.INIT = 16'h8888;
    X_LUT4 C18995(
      .ADR0 (\CRT/ssvga_fifo/N740 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C751/N16 )
    );
    defparam C18985.INIT = 16'h8888;
    X_LUT4 C18985(
      .ADR0 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR1 (\CRT/ssvga_fifo/N741 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C751/N21 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr_plus1<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[3]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<2> (
      .I (\CRT/ssvga_fifo/C751/N16 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [2])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<3> (
      .I (\CRT/ssvga_fifo/C751/N21 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [3])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17657.INIT = 16'h7878;
    X_LUT4 C17657(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [1]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_waddr [0]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_waddr [2]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N306 )
    );
    defparam C17655.INIT = 16'h78F0;
    X_LUT4 C17655(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [1]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_waddr [0]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_waddr [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_waddr [2]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N307 )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/waddr_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N306 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_waddr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr [2])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_waddr<3>/FFY/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[3]/FFY/RST )
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_waddr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_waddr[3]/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/waddr_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N307 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_waddr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr [3])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_waddr<3>/FFX/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[3]/FFX/RST )
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_waddr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_waddr[3]/FFX/RST ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18997.INIT = 16'h8888;
    X_LUT4 C18997(
      .ADR0 (\CRT/ssvga_fifo/N742 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C751/N26 )
    );
    defparam C18983.INIT = 16'hCC00;
    X_LUT4 C18983(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/N743 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .O (\CRT/ssvga_fifo/C751/N31 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr_plus1<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[5]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<4> (
      .I (\CRT/ssvga_fifo/C751/N26 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [4])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<5> (
      .I (\CRT/ssvga_fifo/C751/N31 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [5])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17654.INIT = 16'h5AF0;
    X_LUT4 C17654(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [3]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_waddr [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/C332/C3/C1 ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N308 )
    );
    defparam C17656.INIT = 16'h8080;
    X_LUT4 C17656(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_waddr [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_waddr [0]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[4]/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_waddr<4>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_waddr[4]/FROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/C332/C3/C1 )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/waddr_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N308 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_waddr[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr [4])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_waddr<4>/FFY/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[4]/FFY/RST )
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_waddr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_waddr[4]/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17731.INIT = 16'h0FF0;
    X_LUT4 C17731(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [0]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [1]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/GROM )
    );
    defparam \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<0>/F .INIT = 16'h0000;
    X_LUT4 \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<0>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<0>/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/GROM ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next [0])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FROM ),
      .O (GLOBAL_LOGIC0_7)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/waddr_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18996.INIT = 16'hAA00;
    X_LUT4 C18996(
      .ADR0 (\CRT/ssvga_fifo/N744 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .O (\CRT/ssvga_fifo/C751/N36 )
    );
    defparam C18984.INIT = 16'h8888;
    X_LUT4 C18984(
      .ADR0 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR1 (\CRT/ssvga_fifo/N745 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C751/N41 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr_plus1<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[7]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<6> (
      .I (\CRT/ssvga_fifo/C751/N36 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [6])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<7> (
      .I (\CRT/ssvga_fifo/C751/N41 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [7])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17729.INIT = 16'h5FA0;
    X_LUT4 C17729(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [0]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [1]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [2]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N288 )
    );
    defparam C17727.INIT = 16'h6AAA;
    X_LUT4 C17727(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [3]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [1]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [0]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [2]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N289 )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_waddr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/waddr_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N288 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr [2])
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbw_waddr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/waddr_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N289 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/FFX/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr [3])
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbw_waddr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18224.INIT = 16'h0010;
    X_LUT4 C18224(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [7]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [6]),
      .ADR2 (syn181347),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 ),
      .O (N12588)
    );
    defparam C18226.INIT = 16'h0055;
    X_LUT4 C18226(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/S_19/cell0 )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out_reg (
      .I (N12588),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/FFY/ASYNC_FF_GSR_OR_25 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C18982.INIT = 16'h8888;
    X_LUT4 C18982(
      .ADR0 (\CRT/ssvga_fifo/N746 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C751/N46 )
    );
    defparam C19000.INIT = 16'hCC00;
    X_LUT4 C19000(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/N747 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .O (\CRT/ssvga_fifo/C751/N51 )
    );
    X_INV \CRT/ssvga_fifo/rd_ptr_plus1<9>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[9]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<8> (
      .I (\CRT/ssvga_fifo/C751/N46 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [8])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/rd_ptr_plus1_reg<9> (
      .I (\CRT/ssvga_fifo/C751/N51 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12082),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ptr_plus1[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1 [9])
    );
    X_OR2 \CRT/ssvga_fifo/rd_ptr_plus1<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/rd_ptr_plus1[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17726.INIT = 16'h3CF0;
    X_LUT4 C17726(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [4]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/C310/C3/C1 ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N290 )
    );
    defparam C17728.INIT = 16'hA000;
    X_LUT4 C17728(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [0]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [1]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_waddr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_waddr<4>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/C310/C3/C1 )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/waddr_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N290 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr [4])
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbw_waddr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18268.INIT = 16'hFFA0;
    X_LUT4 C18268(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/C14/N24 ),
      .ADR3 (syn181285),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/GROM )
    );
    defparam C18269.INIT = 16'h0C0A;
    X_LUT4 C18269(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be [0]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [0]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (syn18908),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_be_out<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_be_out<0>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_be_out [0])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_be_out<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/FROM ),
      .O (syn181285)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/be_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out [0])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_be_out<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17635.INIT = 16'h2222;
    X_LUT4 C17635(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wclock_nempty_detect )
      ,
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty121 )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty_reg (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty121 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR_26 (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C18263.INIT = 16'hFF88;
    X_LUT4 C18263(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/C14/N18 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR2 (VCC),
      .ADR3 (syn181298),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/GROM )
    );
    defparam C18264.INIT = 16'h0E04;
    X_LUT4 C18264(
      .ADR0 (syn18908),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be [1]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [1]),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_be_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_be_out<1>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_be_out [1])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_be_out<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/FROM ),
      .O (syn181298)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/be_out_reg<1> (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out [1])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_be_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18258.INIT = 16'hFFC0;
    X_LUT4 C18258(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/C14/N12 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (syn181311),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/GROM )
    );
    defparam C18259.INIT = 16'h0A0C;
    X_LUT4 C18259(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [2]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be [2]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (syn18908),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_be_out<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_be_out<2>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_be_out [2])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_be_out<2>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/FROM ),
      .O (syn181311)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/be_out_reg<2> (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out [2])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_be_out<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[2]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17901.INIT = 16'hFFC0;
    X_LUT4 C17901(
      .ADR0 (VCC),
      .ADR1 (syn22790),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR3 (syn182097),
      .O (\bridge/pci_target_unit/wishbone_master/C83/N38 )
    );
    defparam C17902.INIT = 16'hFCF8;
    X_LUT4 C17902(
      .ADR0 (syn17020),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C983 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .ADR3 (syn17011),
      .O (\bridge/pci_target_unit/wishbone_master/c_state[0]/FROM )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/c_state<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/c_state[0]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/c_state<0>/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/c_state[0]/FROM ),
      .O (syn182097)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/c_state_reg<0> (
      .I (\bridge/pci_target_unit/wishbone_master/C83/N38 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/c_state[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/c_state [0])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/c_state<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/c_state[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/c_state[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18253.INIT = 16'hFFC0;
    X_LUT4 C18253(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/C14/N6 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (syn181324),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/GROM )
    );
    defparam C18254.INIT = 16'h5044;
    X_LUT4 C18254(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [3]),
      .ADR3 (syn18908),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_be_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_be_out<3>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_be_out [3])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_be_out<3>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/FROM ),
      .O (syn181324)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/be_out_reg<3> (
      .I (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out [3])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_be_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_be_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17897.INIT = 16'hFFE0;
    X_LUT4 C17897(
      .ADR0 (\bridge/pci_target_unit/del_sync_bc_out [0]),
      .ADR1 (syn19710),
      .ADR2 (syn17090),
      .ADR3 (syn182109),
      .O (\bridge/pci_target_unit/wishbone_master/C83/N27 )
    );
    defparam C17898.INIT = 16'hFEEE;
    X_LUT4 C17898(
      .ADR0 (syn182107),
      .ADR1 (syn22805),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C983 ),
      .ADR3 (syn17020),
      .O (\bridge/pci_target_unit/wishbone_master/c_state[1]/FROM )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/c_state<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/c_state[1]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/c_state<1>/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/c_state[1]/FROM ),
      .O (syn182109)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/c_state_reg<1> (
      .I (\bridge/pci_target_unit/wishbone_master/C83/N27 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/c_state[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/c_state [1])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/c_state<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/c_state[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/c_state[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17906.INIT = 16'hEAAA;
    X_LUT4 C17906(
      .ADR0 (syn22771),
      .ADR1 (syn19580),
      .ADR2 (\bridge/pci_target_unit/del_sync_comp_req_pending_out ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/c_state [2]),
      .O (\bridge/pci_target_unit/wishbone_master/C83/N15 )
    );
    defparam C19255.INIT = 16'h0050;
    X_LUT4 C19255(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/c_state [0]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/c_state [1]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/c_state [2]),
      .O (\bridge/pci_target_unit/wishbone_master/c_state[2]/FROM )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/c_state<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/c_state[2]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/c_state<2>/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/c_state[2]/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C977 )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/c_state_reg<2> (
      .I (\bridge/pci_target_unit/wishbone_master/C83/N15 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/c_state[2]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/c_state [2])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/c_state<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/c_state[2]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/c_state[2]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18202.INIT = 16'h33CC;
    X_LUT4 C18202(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [0]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/GROM )
    );
    defparam \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<1>/F .INIT = 16'h0000;
    X_LUT4 \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<1>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<1>/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/GROM ),
      .O (\bridge/wishbone_slave_unit/fifos/inNextGreyCount [0])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FROM ),
      .O (GLOBAL_LOGIC0_11)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/inGreyCount_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/in_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/inNextGreyCount [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/in_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18194.INIT = 16'h0FF0;
    X_LUT4 C18194(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [1]),
      .O (\bridge/wishbone_slave_unit/fifos/inNextGreyCount [1])
    );
    X_INV \bridge/wishbone_slave_unit/fifos/inGreyCount<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/inGreyCount_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/inNextGreyCount [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/in_count_en ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/inGreyCount[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount [1])
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/inGreyCount<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/inGreyCount[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18204.INIT = 16'h5A5A;
    X_LUT4 C18204(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [3]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/inNextGreyCount [2])
    );
    X_INV \bridge/wishbone_slave_unit/fifos/inGreyCount<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/inGreyCount_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/inNextGreyCount [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/in_count_en ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/inGreyCount[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount [2])
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/inGreyCount<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/inGreyCount[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/inGreyCount_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/in_count_en ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/inGreyCount[3]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount [3])
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/inGreyCount<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/inGreyCount[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/inGreyCount[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18839.INIT = 16'hA0A0;
    X_LUT4 C18839(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (VCC),
      .O (\bridge/configuration/C384/N3 )
    );
    defparam C18823.INIT = 16'hF000;
    X_LUT4 C18823(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .O (\bridge/configuration/C383/N3 )
    );
    X_INV \bridge/configuration/delete_status_bit13/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/delete_status_bit13/SRNOT )
    );
    X_FF \bridge/configuration/delete_status_bit12_reg (
      .I (\bridge/configuration/C384/N3 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C338/N3 ),
      .SET (\bridge/configuration/delete_status_bit13/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_status_bit12 )
    );
    X_OR2 \bridge/configuration/delete_status_bit13/FFY/ASYNC_FF_GSR_OR_27 (
      .I0 (\bridge/configuration/delete_status_bit13/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_status_bit13/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/delete_status_bit13_reg (
      .I (\bridge/configuration/C383/N3 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C338/N3 ),
      .SET (\bridge/configuration/delete_status_bit13/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_status_bit13 )
    );
    X_OR2 \bridge/configuration/delete_status_bit13/FFX/ASYNC_FF_GSR_OR_28 (
      .I0 (\bridge/configuration/delete_status_bit13/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_status_bit13/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18135.INIT = 16'h0101;
    X_LUT4 C18135(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/lock ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending ),
      .ADR3 (VCC),
      .O (N12589)
    );
    defparam C18138.INIT = 16'h1000;
    X_LUT4 C18138(
      .ADR0 (syn19577),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending ),
      .ADR3 (syn17678),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/wdel_completion_allow )
    );
    X_INV
     \bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/do_del_request_reg (
      .I (N12589),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/wishbone_slave/do_del_request )
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/FFY/ASYNC_FF_GSR_OR_29 (
      .I0 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow_reg (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/wdel_completion_allow ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow )
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/FFX/ASYNC_FF_GSR_OR_30 (
      .I0 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow/FFX/ASYNC_FF_GSR_OR )

    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_sm/ad_iob_oe_feed/C40 .INIT = 16'hFF80;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_sm/ad_iob_oe_feed/C40 (
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep ),
      .ADR1 (N_STOP),
      .ADR2 (N_TRDY),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_slow ),
      .O (\bridge/output_backup/mas_ad_en_out/GROM )
    );
    defparam C19453.INIT = 16'hFFF8;
    X_LUT4 C19453(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_bc_out [0]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C4/N9 ),
      .ADR2 (syn18939),
      .ADR3 (syn18937),
      .O (\bridge/output_backup/mas_ad_en_out/FROM )
    );
    X_INV \bridge/output_backup/mas_ad_en_out/SRMUX (
      .I (N_RST),
      .O (\bridge/output_backup/mas_ad_en_out/SRNOT )
    );
    X_BUF \bridge/output_backup/mas_ad_en_out/YUSED (
      .I (\bridge/output_backup/mas_ad_en_out/GROM ),
      .O (\bridge/pci_mux_mas_ad_en_in )
    );
    X_BUF \bridge/output_backup/mas_ad_en_out/XUSED (
      .I (\bridge/output_backup/mas_ad_en_out/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_slow )
    );
    X_FF \bridge/output_backup/mas_ad_en_out_reg (
      .I (\bridge/output_backup/mas_ad_en_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/output_backup/mas_ad_en_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/output_backup/mas_ad_en_out )
    );
    X_OR2 \bridge/output_backup/mas_ad_en_out/FFY/ASYNC_FF_GSR_OR_31 (
      .I0 (\bridge/output_backup/mas_ad_en_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/output_backup/mas_ad_en_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17677.INIT = 16'h5500;
    X_LUT4 C17677(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect )
      ,
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty116 )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty_reg (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty116 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR_32 (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C19035.INIT = 16'hFFAA;
    X_LUT4 C19035(
      .ADR0 (\CRT/ssvga_wbm_if/N1515 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1474/N6 )
    );
    defparam C19051.INIT = 16'hEEEE;
    X_LUT4 C19051(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1516 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N11 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[1]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<0> (
      .I (\CRT/ssvga_wbm_if/C1474/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [0])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<1> (
      .I (\CRT/ssvga_wbm_if/C1474/N11 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[1]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [1])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17742.INIT = 16'hEECC;
    X_LUT4 C17742(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .ADR1 (syn23263),
      .ADR2 (VCC),
      .ADR3 (syn182435),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/reg_full )
    );
    defparam C17743.INIT = 16'h8008;
    X_LUT4 C17743(
      .ADR0 (syn182431),
      .ADR1 (syn182432),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [0]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [0]),
      .O (\bridge/wishbone_slave_unit/fifos_wbw_full_out/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/fifos_wbw_full_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos_wbw_full_out/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos_wbw_full_out/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos_wbw_full_out/FROM ),
      .O (syn182435)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/full_reg (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/reg_full ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos_wbw_full_out/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos_wbw_full_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos_wbw_full_out/FFY/ASYNC_FF_GSR_OR_33 (
      .I0 (\bridge/wishbone_slave_unit/fifos_wbw_full_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos_wbw_full_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19309.INIT = 16'h555D;
    X_LUT4 C19309(
      .ADR0 (syn178884),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .ADR2 (syn19397),
      .ADR3 (syn19385),
      .O (\bridge/pci_target_unit/fifos/pciw_write_performed/GROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_write_performed/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_write_performed/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_write_performed/BYMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_write_performed/BYNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_write_performed/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_write_performed/GROM ),
      .O (N12616)
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_write_performed_reg (
      .I (\bridge/pci_target_unit/fifos/pciw_write_performed/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_write_performed/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_write_performed )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_write_performed/FFY/ASYNC_FF_GSR_OR_34 (
      .I0 (\bridge/pci_target_unit/fifos/pciw_write_performed/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_write_performed/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19031.INIT = 16'hFFAA;
    X_LUT4 C19031(
      .ADR0 (\CRT/ssvga_wbm_if/N1517 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1474/N16 )
    );
    defparam C19055.INIT = 16'hEEEE;
    X_LUT4 C19055(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1518 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N21 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[3]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<2> (
      .I (\CRT/ssvga_wbm_if/C1474/N16 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [2])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<3> (
      .I (\CRT/ssvga_wbm_if/C1474/N21 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[3]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [3])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/serr_en_crit_gen/C32 .INIT = 16'h0AA0;
    X_LUT4 \bridge/parity_checker/serr_en_crit_gen/C32 (
      .ADR0 (\bridge/parity_checker/serr_generate ),
      .ADR1 (VCC),
      .ADR2 (\bridge/parity_checker/non_critical_par ),
      .ADR3 (N_PAR),
      .O (\bridge/parchk_sig_serr_out/GROM )
    );
    X_INV \bridge/parchk_sig_serr_out/SRMUX (
      .I (N_RST),
      .O (\bridge/parchk_sig_serr_out/SRNOT )
    );
    X_BUF \bridge/parchk_sig_serr_out/YUSED (
      .I (\bridge/parchk_sig_serr_out/GROM ),
      .O (\bridge/pci_mux_serr_en_in )
    );
    X_FF \bridge/output_backup/serr_en_out_reg (
      .I (\bridge/parchk_sig_serr_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/parchk_sig_serr_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/parchk_sig_serr_out )
    );
    X_OR2 \bridge/parchk_sig_serr_out/FFY/ASYNC_FF_GSR_OR_35 (
      .I0 (\bridge/parchk_sig_serr_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/parchk_sig_serr_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19033.INIT = 16'hFFAA;
    X_LUT4 C19033(
      .ADR0 (\CRT/ssvga_wbm_if/N1519 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1474/N26 )
    );
    defparam C19052.INIT = 16'hFFCC;
    X_LUT4 C19052(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_wbm_if/N1520 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1474/N31 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[5]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<4> (
      .I (\CRT/ssvga_wbm_if/C1474/N26 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[5]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [4])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<5> (
      .I (\CRT/ssvga_wbm_if/C1474/N31 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[5]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [5])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19157.INIT = 16'h2222;
    X_LUT4 C19157(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/GROM )
    );
    defparam C19320.INIT = 16'h8888;
    X_LUT4 C19320(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/pci_target_sm/N63 )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/state_backoff_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/state_backoff_reg/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/GROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/N64 )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/state_transfere_reg_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/state_transfere_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/state_backoff_reg/FFY/ASYNC_FF_GSR_OR_36 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/state_backoff_reg_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/N63 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/state_backoff_reg/FFX/ASYNC_FF_GSR_OR_37 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_sm/cbe_iob_feed/C40 .INIT = 16'hFF80;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_sm/cbe_iob_feed/C40 (
      .ADR0 (N_STOP),
      .ADR1 (N_TRDY),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/frame_en_keep ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cbe_en_slow ),
      .O (\bridge/out_bckp_cbe_en_out/GROM )
    );
    defparam C19455.INIT = 16'hFFFE;
    X_LUT4 C19455(
      .ADR0 (syn18930),
      .ADR1 (syn18937),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .ADR3 (syn18939),
      .O (\bridge/out_bckp_cbe_en_out/FROM )
    );
    X_INV \bridge/out_bckp_cbe_en_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_cbe_en_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_cbe_en_out/YUSED (
      .I (\bridge/out_bckp_cbe_en_out/GROM ),
      .O (\bridge/pci_mux_cbe_en_in )
    );
    X_BUF \bridge/out_bckp_cbe_en_out/XUSED (
      .I (\bridge/out_bckp_cbe_en_out/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cbe_en_slow )
    );
    X_FF \bridge/output_backup/cbe_en_out_reg (
      .I (\bridge/out_bckp_cbe_en_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/out_bckp_cbe_en_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_cbe_en_out )
    );
    X_OR2 \bridge/out_bckp_cbe_en_out/FFY/ASYNC_FF_GSR_OR_38 (
      .I0 (\bridge/out_bckp_cbe_en_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_cbe_en_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18913.INIT = 16'hAA00;
    X_LUT4 C18913(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .O (\bridge/configuration/C382/N3 )
    );
    defparam C18817.INIT = 16'h8888;
    X_LUT4 C18817(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/configuration/C381/N3 )
    );
    X_INV \bridge/configuration/delete_status_bit15/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/delete_status_bit15/SRNOT )
    );
    X_FF \bridge/configuration/delete_status_bit14_reg (
      .I (\bridge/configuration/C382/N3 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C338/N3 ),
      .SET (\bridge/configuration/delete_status_bit15/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_status_bit14 )
    );
    X_OR2 \bridge/configuration/delete_status_bit15/FFY/ASYNC_FF_GSR_OR_39 (
      .I0 (\bridge/configuration/delete_status_bit15/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_status_bit15/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/delete_status_bit15_reg (
      .I (\bridge/configuration/C381/N3 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C338/N3 ),
      .SET (\bridge/configuration/delete_status_bit15/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_status_bit15 )
    );
    X_OR2 \bridge/configuration/delete_status_bit15/FFX/ASYNC_FF_GSR_OR_40 (
      .I0 (\bridge/configuration/delete_status_bit15/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_status_bit15/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19032.INIT = 16'hFAFA;
    X_LUT4 C19032(
      .ADR0 (\CRT/ssvga_wbm_if/N1521 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N36 )
    );
    defparam C19053.INIT = 16'hFFF0;
    X_LUT4 C19053(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (\CRT/ssvga_wbm_if/N1522 ),
      .O (\CRT/ssvga_wbm_if/C1474/N41 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[7]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<6> (
      .I (\CRT/ssvga_wbm_if/C1474/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[7]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [6])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<7> (
      .I (\CRT/ssvga_wbm_if/C1474/N41 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[7]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [7])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19050.INIT = 16'hFAFA;
    X_LUT4 C19050(
      .ADR0 (\CRT/ssvga_wbm_if/N1523 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N46 )
    );
    defparam C19034.INIT = 16'hEEEE;
    X_LUT4 C19034(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1524 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N51 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<9>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[9]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<8> (
      .I (\CRT/ssvga_wbm_if/C1474/N46 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[9]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [8])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<9> (
      .I (\CRT/ssvga_wbm_if/C1474/N51 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[9]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [9])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18217.INIT = 16'h0500;
    X_LUT4 C18217(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/decode_count [1]),
      .ADR3 (syn17018),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/do_master_abort )
    );
    defparam C18218.INIT = 16'hA000;
    X_LUT4 C18218(
      .ADR0 (N_TRDY),
      .ADR1 (VCC),
      .ADR2 (N_STOP),
      .ADR3 (N_DEVSEL),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FROM ),
      .O (syn17018)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/mabort1_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/do_master_abort ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FFY/ASYNC_FF_GSR_OR_41 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2 )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FFX/ASYNC_FF_GSR_OR_42 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17910.INIT = 16'hDDCD;
    X_LUT4 C17910(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/stop_w ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_89/cell0 ),
      .O (\bridge/pci_target_unit/pci_target_sm/C4/N19 )
    );
    defparam C17911.INIT = 16'hF3F1;
    X_LUT4 C17911(
      .ADR0 (syn24524),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR2 (\bridge/pci_target_unit/pcit_if_disconect_wo_data_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_pcir_fifo_data_err_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/c_state[0]/FROM )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/c_state<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/c_state[0]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/c_state<0>/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/c_state[0]/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/S_89/cell0 )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/c_state_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_sm/C4/N19 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/c_state[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/c_state [0])
    );
    X_OR2 \bridge/pci_target_unit/pci_target_sm/c_state<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_sm/c_state[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pci_target_sm/c_state[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17909.INIT = 16'h22CC;
    X_LUT4 C17909(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_89/cell0 ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .O (\bridge/pci_target_unit/pci_target_sm/C4/N11 )
    );
    defparam C19129.INIT = 16'h0C00;
    X_LUT4 C19129(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR2 (\bridge/out_bckp_stop_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .O (\bridge/pci_target_unit/pci_target_sm/c_state[1]/FROM )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/c_state<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/c_state[1]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/c_state<1>/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/c_state[1]/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/stop_w_frm )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/c_state_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_sm/C4/N11 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/c_state[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/c_state [1])
    );
    X_OR2 \bridge/pci_target_unit/pci_target_sm/c_state<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_sm/c_state[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pci_target_sm/c_state[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17757.INIT = 16'hF333;
    X_LUT4 C17757(
      .ADR0 (VCC),
      .ADR1 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect80 ),
      .ADR2 (syn19088),
      .ADR3 (syn182406),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/reg_empty )
    );
    defparam C18201.INIT = 16'hC0C0;
    X_LUT4 C18201(
      .ADR0 (VCC),
      .ADR1 (syn19088),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_control_out [0]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/out_count_en )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty_reg (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/reg_empty ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR_43 (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19044.INIT = 16'h2222;
    X_LUT4 C19044(
      .ADR0 (\CRT/ssvga_wbm_if/N1525 ),
      .ADR1 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N56 )
    );
    defparam C19048.INIT = 16'hEEEE;
    X_LUT4 C19048(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1526 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N62 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<11>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[11]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<10> (
      .I (\CRT/ssvga_wbm_if/C1474/N56 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST (\CRT/ssvga_wbm_if/vmaddr_r[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [10])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[11]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<11> (
      .I (\CRT/ssvga_wbm_if/C1474/N62 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[11]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [11])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[11]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18021.INIT = 16'hFF80;
    X_LUT4 C18021(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [2]),
      .ADR3 (syn181803),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N6 )
    );
    defparam C18022.INIT = 16'h7340;
    X_LUT4 C18022(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [2]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3384 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[2]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[2]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<2>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[2]/FROM ),
      .O (syn181803)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<2> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[2]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[2]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[2]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18018.INIT = 16'hFF80;
    X_LUT4 C18018(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [3]),
      .ADR3 (syn181810),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N12 )
    );
    defparam C18019.INIT = 16'h4F40;
    X_LUT4 C18019(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [3]),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3385 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[3]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[3]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<3>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[3]/FROM ),
      .O (syn181810)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<3> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19045.INIT = 16'h4444;
    X_LUT4 C19045(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1527 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N66 )
    );
    defparam C19047.INIT = 16'hEEEE;
    X_LUT4 C19047(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1528 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N72 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<13>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[13]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<12> (
      .I (\CRT/ssvga_wbm_if/C1474/N66 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST (\CRT/ssvga_wbm_if/vmaddr_r[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [12])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[13]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<13> (
      .I (\CRT/ssvga_wbm_if/C1474/N72 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[13]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [13])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[13]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[13]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18016.INIT = 16'hFF80;
    X_LUT4 C18016(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [4]),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (syn181815),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N18 )
    );
    defparam C18017.INIT = 16'h30B8;
    X_LUT4 C18017(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [4]),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3386 ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[4]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[4]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<4>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[4]/FROM ),
      .O (syn181815)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<4> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18014.INIT = 16'hFF80;
    X_LUT4 C18014(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [5]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (syn181820),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N24 )
    );
    defparam C18015.INIT = 16'h3A0A;
    X_LUT4 C18015(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3387 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [5]),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[5]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[5]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<5>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[5]/FROM ),
      .O (syn181820)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<5> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N24 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [5])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19036.INIT = 16'h0A0A;
    X_LUT4 C19036(
      .ADR0 (\CRT/ssvga_wbm_if/N1529 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N76 )
    );
    defparam C19049.INIT = 16'h0C0C;
    X_LUT4 C19049(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_wbm_if/N1530 ),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N81 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<15>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[15]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<14> (
      .I (\CRT/ssvga_wbm_if/C1474/N76 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST (\CRT/ssvga_wbm_if/vmaddr_r[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [14])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[15]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<15> (
      .I (\CRT/ssvga_wbm_if/C1474/N81 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST (\CRT/ssvga_wbm_if/vmaddr_r[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [15])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[15]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[15]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17787.INIT = 16'hCCFF;
    X_LUT4 C17787(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/comp_done_reg_clr ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/comp_done_reg_main ),
      .O (N12603)
    );
    defparam C17786.INIT = 16'hDC50;
    X_LUT4 C17786(
      .ADR0 (\bridge/pci_target_unit/del_sync/comp_done_reg_clr ),
      .ADR1 (syn22771),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_done_reg_main ),
      .ADR3 (\bridge/pci_target_unit/del_sync_comp_req_pending_out ),
      .O (\bridge/pciu_pci_drcomp_pending_out/FROM )
    );
    X_INV \bridge/pciu_pci_drcomp_pending_out/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_pci_drcomp_pending_out/SRNOT )
    );
    X_BUF \bridge/pciu_pci_drcomp_pending_out/XUSED (
      .I (\bridge/pciu_pci_drcomp_pending_out/FROM ),
      .O (N12542)
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_comp_pending_reg (
      .I (N12603),
      .CLK (CLK_BUFGPed),
      .CE (N12542),
      .SET (GND),
      .RST (\bridge/pciu_pci_drcomp_pending_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_pci_drcomp_pending_out )
    );
    X_OR2 \bridge/pciu_pci_drcomp_pending_out/FFY/ASYNC_FF_GSR_OR_44 (
      .I0 (\bridge/pciu_pci_drcomp_pending_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_pci_drcomp_pending_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18012.INIT = 16'hFF80;
    X_LUT4 C18012(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [6]),
      .ADR3 (syn181825),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N30 )
    );
    defparam C18013.INIT = 16'h44E4;
    X_LUT4 C18013(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3388 ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [6]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[6]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<6>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[6]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<6>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[6]/FROM ),
      .O (syn181825)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<6> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[6]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [6])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<6>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[6]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[6]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18010.INIT = 16'hFF80;
    X_LUT4 C18010(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [7]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (syn181830),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N36 )
    );
    defparam C18011.INIT = 16'h44F0;
    X_LUT4 C18011(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [7]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3389 ),
      .ADR3 (N12594),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[7]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[7]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<7>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[7]/FROM ),
      .O (syn181830)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<7> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [7])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19046.INIT = 16'hFAFA;
    X_LUT4 C19046(
      .ADR0 (\CRT/ssvga_wbm_if/N1531 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1474/N87 )
    );
    X_INV \CRT/ssvga_wbm_if/vmaddr_r<16>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[16]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/vmaddr_r_reg<16> (
      .I (\CRT/ssvga_wbm_if/C1474/N87 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (\CRT/ssvga_wbm_if/vmaddr_r[16]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_wbm_if/vmaddr_r [16])
    );
    X_OR2 \CRT/ssvga_wbm_if/vmaddr_r<16>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_wbm_if/vmaddr_r[16]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_wbm_if/vmaddr_r[16]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18008.INIT = 16'hFF80;
    X_LUT4 C18008(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [8]),
      .ADR3 (syn181835),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N42 )
    );
    defparam C18009.INIT = 16'h44F0;
    X_LUT4 C18009(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [8]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3390 ),
      .ADR3 (N12594),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[8]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<8>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[8]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<8>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[8]/FROM ),
      .O (syn181835)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<8> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N42 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[8]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [8])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<8>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[8]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[8]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17646.INIT = 16'h5A5A;
    X_LUT4 C17646(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_waddr [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_waddr [1]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next [1])
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<1>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C18006.INIT = 16'hFF80;
    X_LUT4 C18006(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [9]),
      .ADR3 (syn181840),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N48 )
    );
    defparam C18007.INIT = 16'h0ACA;
    X_LUT4 C18007(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3391 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [9]),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[9]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[9]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<9>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[9]/FROM ),
      .O (syn181840)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<9> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N48 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [9])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[9]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17621.INIT = 16'h55AA;
    X_LUT4 C17621(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_waddr [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_waddr [2]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next [2])
    );
    defparam C17642.INIT = 16'h3C3C;
    X_LUT4 C17642(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_waddr [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_waddr [3]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next [3])
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<3>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_wgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19999.INIT = 16'h4040;
    X_LUT4 C19999(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/map ),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en ),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/pref_en ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out[3]/GROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_bc_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out[3]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_bc_out<3>/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_bc_out[3]/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_del_bc_out [3])
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/bc_out_reg<3> (
      .I (\bridge/wishbone_slave_unit/del_sync_bc_out[3]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/del_sync_bc_out[3]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out [3])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_bc_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17789.INIT = 16'h0050;
    X_LUT4 C17789(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/S_198/cell0 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/sync_req_comp_pending ),
      .ADR3 (\bridge/pci_target_unit/del_sync/comp_cycle_count [16]),
      .O (\bridge/pci_target_unit/del_sync/C9/N5 )
    );
    X_INV \bridge/pci_target_unit/del_sync/req_comp_pending/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/req_comp_pending/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/req_comp_pending_reg (
      .I (\bridge/pci_target_unit/del_sync/C9/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (N12541),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/req_comp_pending/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/req_comp_pending )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/req_comp_pending/FFY/ASYNC_FF_GSR_OR_45 (
      .I0 (\bridge/pci_target_unit/del_sync/req_comp_pending/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/req_comp_pending/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18119.INIT = 16'h5000;
    X_LUT4 C18119(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [16]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending ),
      .ADR3 (syn22126),
      .O (\bridge/wishbone_slave_unit/del_sync/C9/N5 )
    );
    defparam C18120.INIT = 16'hAF23;
    X_LUT4 C18120(
      .ADR0 (syn181420),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/C707 ),
      .ADR2 (syn16935),
      .ADR3 (\bridge/wishbone_slave_unit/wishbone_slave/C749 ),
      .O (\bridge/wishbone_slave_unit/del_sync/req_comp_pending/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/req_comp_pending/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/req_comp_pending/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/req_comp_pending/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/req_comp_pending/FROM ),
      .O (syn22126)
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/req_comp_pending_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/C9/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (N12380),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/req_comp_pending/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/req_comp_pending )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/req_comp_pending/FFY/ASYNC_FF_GSR_OR_46 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/req_comp_pending/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17926.INIT = 16'h5F4C;
    X_LUT4 C17926(
      .ADR0 (syn19590),
      .ADR1 (syn182037),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_control_out [0]),
      .ADR3 (syn182038),
      .O (\bridge/pci_target_unit/fifos/C2/N5 )
    );
    defparam C17927.INIT = 16'h7DBE;
    X_LUT4 C17927(
      .ADR0 (\bridge/pci_target_unit/fifos/outGreyCount [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/outGreyCount [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/inGreyCount [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/inGreyCount [0]),
      .O (\bridge/pci_target_unit/del_sync_comp_flush_out/FROM )
    );
    X_INV \bridge/pci_target_unit/del_sync_comp_flush_out/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_comp_flush_out/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/del_sync_comp_flush_out/XUSED (
      .I (\bridge/pci_target_unit/del_sync_comp_flush_out/FROM ),
      .O (syn182038)
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_transaction_ready_out_reg (
      .I (\bridge/pci_target_unit/fifos/C2/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync_comp_flush_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos_pciw_transaction_ready_out )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync_comp_flush_out/FFY/ASYNC_FF_GSR_OR_47 (
      .I0 (\bridge/pci_target_unit/del_sync_comp_flush_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_comp_flush_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_flush_out_reg (
      .I (\bridge/pci_target_unit/del_sync/comp_cycle_count [16]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync_comp_flush_out/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_comp_flush_out )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync_comp_flush_out/FFX/ASYNC_FF_GSR_OR_48 (
      .I0 (\bridge/pci_target_unit/del_sync_comp_flush_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_comp_flush_out/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18181.INIT = 16'h2000;
    X_LUT4 C18181(
      .ADR0 (syn181420),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/C749 ),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/C707 ),
      .ADR3 (syn17678),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C93/N5 )
    );
    X_INV \bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/wbr_fifo_flush_out_reg (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/C93/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out/FFY/ASYNC_FF_GSR_OR_49 (
      .I0 (\bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18189.INIT = 16'h7788;
    X_LUT4 C18189(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [1]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [0]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [2]),
      .O (\bridge/wishbone_slave_unit/fifos/N1860 )
    );
    defparam C18188.INIT = 16'h7F80;
    X_LUT4 C18188(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [1]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [0]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [3]),
      .O (\bridge/wishbone_slave_unit/fifos/N1861 )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/N1860 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/in_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/N1861 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/in_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17623.INIT = 16'hCFCC;
    X_LUT4 C17623(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0 ),
      .ADR2 (N12616),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_95/cell0 ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_almost_full_in )
    );
    defparam C17624.INIT = 16'h8200;
    X_LUT4 C17624(
      .ADR0 (syn182662),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [0]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [0]),
      .ADR3 (syn182663),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_95/cell0 )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_full_reg (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_almost_full_in ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_full )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FFY/ASYNC_FF_GSR_OR_50 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/sync_comp_done ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FFX/ASYNC_FF_GSR_OR_51 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18927.INIT = 16'hF000;
    X_LUT4 C18927(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/N400 ),
      .ADR3 (syn20304),
      .O (\CRT/ssvga_crtc/C531/N5 )
    );
    defparam C18928.INIT = 16'hFFFE;
    X_LUT4 C18928(
      .ADR0 (syn179587),
      .ADR1 (\CRT/ssvga_crtc/hcntr [4]),
      .ADR2 (syn48756),
      .ADR3 (\CRT/ssvga_crtc/hcntr [1]),
      .O (\CRT/ssvga_fifo/sync_ssvga_en/FROM )
    );
    X_INV \CRT/ssvga_fifo/sync_ssvga_en/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/sync_ssvga_en/SRNOT )
    );
    X_BUF \CRT/ssvga_fifo/sync_ssvga_en/XUSED (
      .I (\CRT/ssvga_fifo/sync_ssvga_en/FROM ),
      .O (syn20304)
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<0> (
      .I (\CRT/ssvga_crtc/C531/N5 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_ssvga_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [0])
    );
    X_OR2 \CRT/ssvga_fifo/sync_ssvga_en/FFY/ASYNC_FF_GSR_OR_52 (
      .I0 (\CRT/ssvga_fifo/sync_ssvga_en/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_ssvga_en/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/ssvga_enable_sync/sync_data_out_reg<0> (
      .I (N_LED),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_ssvga_en/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_ssvga_en )
    );
    X_OR2 \CRT/ssvga_fifo/sync_ssvga_en/FFX/ASYNC_FF_GSR_OR_53 (
      .I0 (\CRT/ssvga_fifo/sync_ssvga_en/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_ssvga_en/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18142.INIT = 16'hCC00;
    X_LUT4 C18142(
      .ADR0 (VCC),
      .ADR1 (syn24500),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_wb_mem_io1_out ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/n_859 )
    );
    defparam C18152.INIT = 16'h9933;
    X_LUT4 C18152(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [11]),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [11]),
      .ADR2 (VCC),
      .ADR3 (syn24500),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/map/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/wishbone_slave/map/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/map/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/map/XUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/map/FROM ),
      .O (syn176975)
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/map_reg (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/n_859 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/wishbone_slave/map/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/wishbone_slave/map )
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/map/FFY/ASYNC_FF_GSR_OR_54 (
      .I0 (\bridge/wishbone_slave_unit/wishbone_slave/map/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/map/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18926.INIT = 16'hAA00;
    X_LUT4 C18926(
      .ADR0 (syn20304),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/N401 ),
      .O (\CRT/ssvga_crtc/C531/N10 )
    );
    X_INV \CRT/ssvga_crtc/hcntr<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/hcntr[1]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<1> (
      .I (\CRT/ssvga_crtc/C531/N10 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [1])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18925.INIT = 16'hAA00;
    X_LUT4 C18925(
      .ADR0 (\CRT/ssvga_crtc/N402 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn20304),
      .O (\CRT/ssvga_crtc/C531/N15 )
    );
    defparam C18924.INIT = 16'hCC00;
    X_LUT4 C18924(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/N403 ),
      .ADR2 (VCC),
      .ADR3 (syn20304),
      .O (\CRT/ssvga_crtc/C531/N20 )
    );
    X_INV \CRT/ssvga_crtc/hcntr<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/hcntr[3]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<2> (
      .I (\CRT/ssvga_crtc/C531/N15 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [2])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<3> (
      .I (\CRT/ssvga_crtc/C531/N20 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [3])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18923.INIT = 16'hAA00;
    X_LUT4 C18923(
      .ADR0 (\CRT/ssvga_crtc/N404 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn20304),
      .O (\CRT/ssvga_crtc/C531/N25 )
    );
    defparam C18922.INIT = 16'hCC00;
    X_LUT4 C18922(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/N405 ),
      .ADR2 (VCC),
      .ADR3 (syn20304),
      .O (\CRT/ssvga_crtc/C531/N30 )
    );
    X_INV \CRT/ssvga_crtc/hcntr<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/hcntr[5]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<4> (
      .I (\CRT/ssvga_crtc/C531/N25 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [4])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<5> (
      .I (\CRT/ssvga_crtc/C531/N30 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [5])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18921.INIT = 16'hA0A0;
    X_LUT4 C18921(
      .ADR0 (\CRT/ssvga_crtc/N406 ),
      .ADR1 (VCC),
      .ADR2 (syn20304),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/C531/N35 )
    );
    defparam C18920.INIT = 16'hC0C0;
    X_LUT4 C18920(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/N407 ),
      .ADR2 (syn20304),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/C531/N40 )
    );
    X_INV \CRT/ssvga_crtc/hcntr<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/hcntr[7]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<6> (
      .I (\CRT/ssvga_crtc/C531/N35 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [6])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<7> (
      .I (\CRT/ssvga_crtc/C531/N40 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [7])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18919.INIT = 16'hAA00;
    X_LUT4 C18919(
      .ADR0 (\CRT/ssvga_crtc/N408 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn20304),
      .O (\CRT/ssvga_crtc/C531/N45 )
    );
    defparam C18918.INIT = 16'h8888;
    X_LUT4 C18918(
      .ADR0 (syn20304),
      .ADR1 (\CRT/ssvga_crtc/N409 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/C531/N50 )
    );
    X_INV \CRT/ssvga_crtc/hcntr<9>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/hcntr[9]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<8> (
      .I (\CRT/ssvga_crtc/C531/N45 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [8])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/hcntr_reg<9> (
      .I (\CRT/ssvga_crtc/C531/N50 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/hcntr[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/hcntr [9])
    );
    X_OR2 \CRT/ssvga_crtc/hcntr<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/hcntr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/hcntr[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18270.INIT = 16'h5C5C;
    X_LUT4 C18270(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [0]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [0]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/GROM )
    );
    defparam C18265.INIT = 16'h22EE;
    X_LUT4 C18265(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [1]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [1]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FROM )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<1>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/SRNOT )
    );
    X_BUF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<1>/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/GROM )
      ,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C14/N24 )
    );
    X_BUF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FROM )
      ,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C14/N18 )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be_reg<0> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/GROM )
      ,
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be_reg<1> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FROM )
      ,
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18260.INIT = 16'h7722;
    X_LUT4 C18260(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [2]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [2]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/GROM )
    );
    defparam C18255.INIT = 16'h33F0;
    X_LUT4 C18255(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_cbe_out [3]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FROM )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<3>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/SRNOT )
    );
    X_BUF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<3>/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/GROM )
      ,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C14/N12 )
    );
    X_BUF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<3>/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FROM )
      ,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C14/N6 )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be_reg<2> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/GROM )
      ,
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be_reg<3> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FROM )
      ,
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_be[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_control_enable_critical/C50 .INIT = 16'hFF22;
    X_LUT4
     \bridge/pci_target_unit/pci_target_sm/pci_target_control_enable_critical/C50 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR1 (N_IRDY),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/ctrl_en_w ),
      .O (\bridge/out_bckp_trdy_en_out/GROM )
    );
    defparam C19154.INIT = 16'hFAFE;
    X_LUT4 C19154(
      .ADR0 (syn179261),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR2 (syn17093),
      .ADR3 (\bridge/in_reg_frame_out ),
      .O (\bridge/out_bckp_trdy_en_out/FROM )
    );
    X_INV \bridge/out_bckp_trdy_en_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_trdy_en_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_trdy_en_out/YUSED (
      .I (\bridge/out_bckp_trdy_en_out/GROM ),
      .O (\bridge/pciu_pciif_devsel_en_out )
    );
    X_BUF \bridge/out_bckp_trdy_en_out/XUSED (
      .I (\bridge/out_bckp_trdy_en_out/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/ctrl_en_w )
    );
    X_FF \bridge/output_backup/trdy_en_out_reg (
      .I (\bridge/out_bckp_trdy_en_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/out_bckp_trdy_en_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_trdy_en_out )
    );
    X_OR2 \bridge/out_bckp_trdy_en_out/FFY/ASYNC_FF_GSR_OR_55 (
      .I0 (\bridge/out_bckp_trdy_en_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_trdy_en_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19022.INIT = 16'hEE44;
    X_LUT4 C19022(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1725 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/pix_start_addr [10]),
      .O (\CRT/ssvga_wbm_if/C1475/N54 )
    );
    defparam C19021.INIT = 16'hE2E2;
    X_LUT4 C19021(
      .ADR0 (\CRT/ssvga_wbm_if/N1726 ),
      .ADR1 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR2 (\CRT/pix_start_addr [11]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1475/N60 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<10> (
      .I (\CRT/ssvga_wbm_if/C1475/N54 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [10])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<11> (
      .I (\CRT/ssvga_wbm_if/C1475/N60 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [11])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19012.INIT = 16'hCACA;
    X_LUT4 C19012(
      .ADR0 (\CRT/ssvga_wbm_if/N1735 ),
      .ADR1 (\CRT/pix_start_addr [20]),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1475/N114 )
    );
    defparam C19011.INIT = 16'hAACC;
    X_LUT4 C19011(
      .ADR0 (\CRT/pix_start_addr [21]),
      .ADR1 (\CRT/ssvga_wbm_if/N1736 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N120 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<20> (
      .I (\CRT/ssvga_wbm_if/C1475/N114 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [20])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<21> (
      .I (\CRT/ssvga_wbm_if/C1475/N120 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [21])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[21]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19020.INIT = 16'hFC30;
    X_LUT4 C19020(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR2 (\CRT/ssvga_wbm_if/N1727 ),
      .ADR3 (\CRT/pix_start_addr [12]),
      .O (\CRT/ssvga_wbm_if/C1475/N66 )
    );
    defparam C19019.INIT = 16'hEE44;
    X_LUT4 C19019(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1728 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/pix_start_addr [13]),
      .O (\CRT/ssvga_wbm_if/C1475/N72 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<12> (
      .I (\CRT/ssvga_wbm_if/C1475/N66 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [12])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<13> (
      .I (\CRT/ssvga_wbm_if/C1475/N72 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [13])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[13]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/cbe_par_calc/C64 .INIT = 16'hF3C0;
    X_LUT4 \bridge/parity_checker/cbe_par_calc/C64 (
      .ADR0 (VCC),
      .ADR1 (\bridge/out_bckp_cbe_en_out ),
      .ADR2 (\bridge/parity_checker/par_cbe_out ),
      .ADR3 (\bridge/parity_checker/cbe_par_calc/syn118 ),
      .O (\bridge/parity_checker/par_cbe_include )
    );
    defparam \bridge/parity_checker/cbe_par_calc/C65 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/cbe_par_calc/C65 (
      .ADR0 (N_CBE[0]),
      .ADR1 (N_CBE[2]),
      .ADR2 (N_CBE[1]),
      .ADR3 (N_CBE[3]),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FROM ),
      .O (\bridge/parity_checker/cbe_par_calc/syn118 )
    );
    X_FF \bridge/parity_checker/cbe_par_reg_reg (
      .I (\bridge/parity_checker/par_cbe_include ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/parity_checker/cbe_par_reg )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FFY/ASYNC_FF_GSR_OR_56 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FFX/ASYNC_FF_GSR_OR_57 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19002.INIT = 16'hCACA;
    X_LUT4 C19002(
      .ADR0 (\CRT/ssvga_wbm_if/N1745 ),
      .ADR1 (\CRT/pix_start_addr [30]),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1475/N174 )
    );
    defparam C19001.INIT = 16'hDD88;
    X_LUT4 C19001(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/pix_start_addr [31]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/N1746 ),
      .O (\CRT/ssvga_wbm_if/C1475/N180 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<30> (
      .I (\CRT/ssvga_wbm_if/C1475/N174 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [30])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<31> (
      .I (\CRT/ssvga_wbm_if/C1475/N180 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [31])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19010.INIT = 16'hF0AA;
    X_LUT4 C19010(
      .ADR0 (\CRT/ssvga_wbm_if/N1737 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [22]),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N126 )
    );
    defparam C19009.INIT = 16'hAACC;
    X_LUT4 C19009(
      .ADR0 (\CRT/pix_start_addr [23]),
      .ADR1 (\CRT/ssvga_wbm_if/N1738 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N132 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<22> (
      .I (\CRT/ssvga_wbm_if/C1475/N126 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [22])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<23> (
      .I (\CRT/ssvga_wbm_if/C1475/N132 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [23])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[23]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19018.INIT = 16'hF0AA;
    X_LUT4 C19018(
      .ADR0 (\CRT/ssvga_wbm_if/N1729 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [14]),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N78 )
    );
    defparam C19017.INIT = 16'hEE44;
    X_LUT4 C19017(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1730 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/pix_start_addr [15]),
      .O (\CRT/ssvga_wbm_if/C1475/N84 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<14> (
      .I (\CRT/ssvga_wbm_if/C1475/N78 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [14])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<15> (
      .I (\CRT/ssvga_wbm_if/C1475/N84 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [15])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[15]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19008.INIT = 16'hF0AA;
    X_LUT4 C19008(
      .ADR0 (\CRT/ssvga_wbm_if/N1739 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [24]),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N138 )
    );
    defparam C19007.INIT = 16'hAACC;
    X_LUT4 C19007(
      .ADR0 (\CRT/pix_start_addr [25]),
      .ADR1 (\CRT/ssvga_wbm_if/N1740 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N144 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<24> (
      .I (\CRT/ssvga_wbm_if/C1475/N138 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [24])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<25> (
      .I (\CRT/ssvga_wbm_if/C1475/N144 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [25])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[25]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19016.INIT = 16'hFC0C;
    X_LUT4 C19016(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_wbm_if/N1731 ),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (\CRT/pix_start_addr [16]),
      .O (\CRT/ssvga_wbm_if/C1475/N90 )
    );
    defparam C19015.INIT = 16'hCFC0;
    X_LUT4 C19015(
      .ADR0 (VCC),
      .ADR1 (\CRT/pix_start_addr [17]),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (\CRT/ssvga_wbm_if/N1732 ),
      .O (\CRT/ssvga_wbm_if/C1475/N96 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<16> (
      .I (\CRT/ssvga_wbm_if/C1475/N90 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [16])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<17> (
      .I (\CRT/ssvga_wbm_if/C1475/N96 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [17])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[17]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19006.INIT = 16'hAAF0;
    X_LUT4 C19006(
      .ADR0 (\CRT/pix_start_addr [26]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_wbm_if/N1741 ),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N150 )
    );
    defparam C19005.INIT = 16'hCCF0;
    X_LUT4 C19005(
      .ADR0 (VCC),
      .ADR1 (\CRT/pix_start_addr [27]),
      .ADR2 (\CRT/ssvga_wbm_if/N1742 ),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N156 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<26> (
      .I (\CRT/ssvga_wbm_if/C1475/N150 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [26])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<27> (
      .I (\CRT/ssvga_wbm_if/C1475/N156 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [27])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[27]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19014.INIT = 16'hEE22;
    X_LUT4 C19014(
      .ADR0 (\CRT/ssvga_wbm_if/N1733 ),
      .ADR1 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR2 (VCC),
      .ADR3 (\CRT/pix_start_addr [18]),
      .O (\CRT/ssvga_wbm_if/C1475/N102 )
    );
    defparam C19013.INIT = 16'hAACC;
    X_LUT4 C19013(
      .ADR0 (\CRT/pix_start_addr [19]),
      .ADR1 (\CRT/ssvga_wbm_if/N1734 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\CRT/ssvga_wbm_if/C1475/N108 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<18> (
      .I (\CRT/ssvga_wbm_if/C1475/N102 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [18])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<19> (
      .I (\CRT/ssvga_wbm_if/C1475/N108 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [19])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[19]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19004.INIT = 16'hCACA;
    X_LUT4 C19004(
      .ADR0 (\CRT/ssvga_wbm_if/N1743 ),
      .ADR1 (\CRT/pix_start_addr [28]),
      .ADR2 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1475/N162 )
    );
    defparam C19003.INIT = 16'hE4E4;
    X_LUT4 C19003(
      .ADR0 (\CRT/ssvga_wbm_if/frame_read ),
      .ADR1 (\CRT/ssvga_wbm_if/N1744 ),
      .ADR2 (\CRT/pix_start_addr [29]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/C1475/N168 )
    );
    X_INV \bridge/wishbone_slave_unit/wb_addr_dec/addr1<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/SRNOT )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<28> (
      .I (\CRT/ssvga_wbm_if/C1475/N162 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [28])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbm_if/wbm_adr_reg<29> (
      .I (\CRT/ssvga_wbm_if/C1475/N168 ),
      .CLK (CLK_BUFGPed),
      .CE (N12065),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [29])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wb_addr_dec/addr1<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[29]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18089.INIT = 16'h0010;
    X_LUT4 C18089(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/err_recovery ),
      .ADR1 (\bridge/conf_wb_err_pending_out ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out ),
      .ADR3 (syn19075),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/GROM )
    );
    defparam C18659.INIT = 16'h8000;
    X_LUT4 C18659(
      .ADR0 (\bridge/conf_wb_err_pending_out ),
      .ADR1 (syn60038),
      .ADR2 (syn17017),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/data_source/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/data_source/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/GROM ),
      .O (N12426)
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/data_source/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/FROM ),
      .O (syn20738)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_source_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12594),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/data_source )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/data_source/FFY/ASYNC_FF_GSR_OR_58 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/data_source/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18081.INIT = 16'hCE0A;
    X_LUT4 C18081(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/err_recovery ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/S_176/cell0 ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_control_out [0]),
      .ADR3 (syn181630),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C8/N6 )
    );
    defparam C18082.INIT = 16'h0011;
    X_LUT4 C18082(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_last_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last ),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/err_recovery ),
      .O (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/FROM )
    );
    X_INV \bridge/pci_target_unit/del_sync/req_comp_pending_sample/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/del_sync/req_comp_pending_sample/XUSED (
      .I (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/FROM ),
      .O (syn181630)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/err_recovery_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C8/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/err_recovery )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/req_comp_pending_sample/FFY/ASYNC_FF_GSR_OR_59 (
      .I0 (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/req_comp_pending_sample_reg (
      .I (\bridge/pci_target_unit/del_sync/sync_req_comp_pending ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/req_comp_pending_sample )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/req_comp_pending_sample/FFX/ASYNC_FF_GSR_OR_60 (
      .I0 (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/req_comp_pending_sample/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/C1122 .INIT = 16'h0F00;
    X_LUT4 \bridge/parity_checker/C1122 (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (N_PERR),
      .ADR3 (\bridge/parity_checker/check_perr ),
      .O (\bridge/parity_checker/perr_sampled_in )
    );
    X_INV \bridge/parity_checker/perr_sampled/SRMUX (
      .I (N_RST),
      .O (\bridge/parity_checker/perr_sampled/SRNOT )
    );
    X_FF \bridge/parity_checker/perr_sampled_reg (
      .I (\bridge/parity_checker/perr_sampled_in ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/parity_checker/perr_sampled/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/parity_checker/perr_sampled )
    );
    X_OR2 \bridge/parity_checker/perr_sampled/FFY/ASYNC_FF_GSR_OR_61 (
      .I0 (\bridge/parity_checker/perr_sampled/SRNOT ),
      .I1 (GSR),
      .O (\bridge/parity_checker/perr_sampled/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18860.INIT = 16'hA0A0;
    X_LUT4 C18860(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (VCC),
      .O (\bridge/configuration/C386/N3 )
    );
    defparam C18815.INIT = 16'hF000;
    X_LUT4 C18815(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .O (\bridge/configuration/C385/N3 )
    );
    X_INV \bridge/configuration/delete_status_bit11/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/delete_status_bit11/SRNOT )
    );
    X_FF \bridge/configuration/delete_status_bit8_reg (
      .I (\bridge/configuration/C386/N3 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C338/N3 ),
      .SET (\bridge/configuration/delete_status_bit11/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_status_bit8 )
    );
    X_OR2 \bridge/configuration/delete_status_bit11/FFY/ASYNC_FF_GSR_OR_62 (
      .I0 (\bridge/configuration/delete_status_bit11/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_status_bit11/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/delete_status_bit11_reg (
      .I (\bridge/configuration/C385/N3 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C338/N3 ),
      .SET (\bridge/configuration/delete_status_bit11/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_status_bit11 )
    );
    X_OR2 \bridge/configuration/delete_status_bit11/FFX/ASYNC_FF_GSR_OR_63 (
      .I0 (\bridge/configuration/delete_status_bit11/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_status_bit11/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17648.INIT = 16'hFFDE;
    X_LUT4 C17648(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [0]),
      .ADR1 (syn182601),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [0]),
      .ADR3 (syn182602),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/GROM )
    );
    defparam C17647.INIT = 16'h8F8F;
    X_LUT4 C17647(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0 ),
      .ADR2 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wclock_nempty_detect90 ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_empty )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/GROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wclock_nempty_detect90 )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wclock_nempty_detect_reg (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wclock_nempty_detect )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR_64 (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty_reg (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_empty ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/FFX/ASYNC_FF_GSR_OR_65 (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17689.INIT = 16'hFFF6;
    X_LUT4 C17689(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [0]),
      .ADR2 (syn182526),
      .ADR3 (syn182527),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/GROM )
    );
    defparam C17690.INIT = 16'h7BDE;
    X_LUT4 C17690(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [1]),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/FROM )
    );
    X_INV
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/SRNOT )
    );
    X_BUF
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/YUSED (
      .I 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/GROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect85 )
    );
    X_BUF
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/XUSED (
      .I 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/FROM ),
      .O (syn182527)
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect_reg (
      .I 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR_66 (
      .I0 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17721.INIT = 16'hFFFC;
    X_LUT4 C17721(
      .ADR0 (VCC),
      .ADR1 (syn182474),
      .ADR2 (syn182473),
      .ADR3 (syn182475),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/GROM )
    );
    defparam C17722.INIT = 16'h7DBE;
    X_LUT4 C17722(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [0]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [1]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [1]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [0]),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/FROM )
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/SRNOT )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/YUSED (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/GROM ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect70 )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/XUSED (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/FROM ),
      .O (syn182475)
    );
    X_FF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect_reg (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR_67 (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17761.INIT = 16'hFFF6;
    X_LUT4 C17761(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [0]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [0]),
      .ADR2 (syn182394),
      .ADR3 (syn182395),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/GROM )
    );
    defparam C17762.INIT = 16'h7DBE;
    X_LUT4 C17762(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [1]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [1]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [2]),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/FROM )
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/SRNOT )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/YUSED (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/GROM ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect80 )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/XUSED (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/FROM ),
      .O (syn182395)
    );
    X_FF
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect_reg (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR_68 (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C18192.INIT = 16'h5AF0;
    X_LUT4 C18192(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [1]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [0]),
      .O (\bridge/wishbone_slave_unit/fifos/N1828 )
    );
    defparam C18191.INIT = 16'h6CCC;
    X_LUT4 C18191(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [1]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [0]),
      .O (\bridge/wishbone_slave_unit/fifos/N1829 )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/N1828 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/N1829 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17614.INIT = 16'hAFAA;
    X_LUT4 C17614(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_95/cell0 ),
      .ADR1 (VCC),
      .ADR2 (N12616),
      .ADR3 (syn182682),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_two_left_in )
    );
    defparam C17615.INIT = 16'h9000;
    X_LUT4 C17615(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [0]),
      .ADR2 (syn182680),
      .ADR3 (syn182679),
      .O (\bridge/pci_target_unit/fifos_pciw_two_left_out/FROM )
    );
    X_INV \bridge/pci_target_unit/fifos_pciw_two_left_out/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos_pciw_two_left_out/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos_pciw_two_left_out/XUSED (
      .I (\bridge/pci_target_unit/fifos_pciw_two_left_out/FROM ),
      .O (syn182682)
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/two_left_out_reg (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_two_left_in ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos_pciw_two_left_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos_pciw_two_left_out )
    );
    X_OR2
     \bridge/pci_target_unit/fifos_pciw_two_left_out/FFY/ASYNC_FF_GSR_OR_69 (
      .I0 (\bridge/pci_target_unit/fifos_pciw_two_left_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos_pciw_two_left_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18949.INIT = 16'hF0FF;
    X_LUT4 C18949(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn16988),
      .ADR3 (syn16982),
      .O (N12150)
    );
    defparam C18950.INIT = 16'h0008;
    X_LUT4 C18950(
      .ADR0 (\CRT/ssvga_crtc/vcntr [0]),
      .ADR1 (syn16986),
      .ADR2 (\CRT/ssvga_crtc/vcntr [2]),
      .ADR3 (\CRT/ssvga_crtc/vcntr [3]),
      .O (\CRT/crtc_vblank/FROM )
    );
    X_INV \CRT/crtc_vblank/SRMUX (
      .I (N_RST),
      .O (\CRT/crtc_vblank/SRNOT )
    );
    X_BUF \CRT/crtc_vblank/XUSED (
      .I (\CRT/crtc_vblank/FROM ),
      .O (syn16982)
    );
    X_FF \CRT/ssvga_crtc/vblank_reg (
      .I (N12150),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12162),
      .SET (GND),
      .RST (\CRT/crtc_vblank/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/crtc_vblank )
    );
    X_OR2 \CRT/crtc_vblank/FFY/ASYNC_FF_GSR_OR_70 (
      .I0 (\CRT/crtc_vblank/SRNOT ),
      .I1 (GSR),
      .O (\CRT/crtc_vblank/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17637.INIT = 16'h0FF0;
    X_LUT4 C17637(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [0]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [1]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next [0])
    );
    defparam C17622.INIT = 16'h33CC;
    X_LUT4 C17622(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [2]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [1]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next [1])
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17706.INIT = 16'h5500;
    X_LUT4 C17706(
      .ADR0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wclock_nempty_detect ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty101 )
    );
    defparam C19978.INIT = 16'h0303;
    X_LUT4 C19978(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty/FROM )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty/FROM )
      ,
      .O (syn17678)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty_reg (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty101 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR_71 (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17636.INIT = 16'h55AA;
    X_LUT4 C17636(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [2]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next [2])
    );
    defparam C17627.INIT = 16'h55AA;
    X_LUT4 C17627(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [3]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next [3])
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/calc_rgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17929.INIT = 16'h3C3C;
    X_LUT4 C17929(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [2]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/inNextGreyCount [1])
    );
    X_INV \bridge/pci_target_unit/fifos/inGreyCount<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/inGreyCount_reg<1> (
      .I (\bridge/pci_target_unit/fifos/inNextGreyCount [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/in_count_en ),
      .SET (\bridge/pci_target_unit/fifos/inGreyCount[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/inGreyCount [1])
    );
    X_OR2 \bridge/pci_target_unit/fifos/inGreyCount<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/inGreyCount[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17638.INIT = 16'hFAAA;
    X_LUT4 C17638(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .ADR3 (syn182630),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_almost_empty )
    );
    defparam C17639.INIT = 16'h8040;
    X_LUT4 C17639(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [0]),
      .ADR1 (syn182627),
      .ADR2 (syn182628),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/FROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/XUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/FROM ),
      .O (syn182630)
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty_reg (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/reg_almost_empty ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/FFY/ASYNC_FF_GSR_OR_72 (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17936.INIT = 16'h3C3C;
    X_LUT4 C17936(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [3]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/inNextGreyCount [2])
    );
    X_INV \bridge/pci_target_unit/fifos/inGreyCount<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/inGreyCount_reg<2> (
      .I (\bridge/pci_target_unit/fifos/inNextGreyCount [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/in_count_en ),
      .SET (\bridge/pci_target_unit/fifos/inGreyCount[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/inGreyCount [2])
    );
    X_OR2 \bridge/pci_target_unit/fifos/inGreyCount<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/inGreyCount[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/inGreyCount_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/in_count_en ),
      .SET (\bridge/pci_target_unit/fifos/inGreyCount[3]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/inGreyCount [3])
    );
    X_OR2 \bridge/pci_target_unit/fifos/inGreyCount<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/inGreyCount[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/inGreyCount[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_sm/frame_iob_feed/C34 .INIT = 16'h2323;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_sm/frame_iob_feed/C34 (
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame ),
      .ADR1 (N12359),
      .ADR2 (N_STOP),
      .ADR3 (VCC),
      .O (\bridge/out_bckp_frame_out/GROM )
    );
    defparam C18230.INIT = 16'hCFCF;
    X_LUT4 C18230(
      .ADR0 (VCC),
      .ADR1 (N12594),
      .ADR2 (N12359),
      .ADR3 (VCC),
      .O (\bridge/out_bckp_frame_out/FROM )
    );
    X_INV \bridge/out_bckp_frame_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_frame_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_frame_out/YUSED (
      .I (\bridge/out_bckp_frame_out/GROM ),
      .O (\bridge/pci_mux_frame_in )
    );
    X_BUF \bridge/out_bckp_frame_out/XUSED (
      .I (\bridge/out_bckp_frame_out/FROM ),
      .O (N12587)
    );
    X_FF \bridge/output_backup/frame_out_reg (
      .I (\bridge/out_bckp_frame_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_frame_load_in ),
      .SET (\bridge/out_bckp_frame_out/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_frame_out )
    );
    X_OR2 \bridge/out_bckp_frame_out/FFY/ASYNC_FF_GSR_OR_73 (
      .I0 (\bridge/out_bckp_frame_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_frame_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17931.INIT = 16'h0FF0;
    X_LUT4 C17931(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/GROM )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_outTransactionCount<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_outTransactionCount<1>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/GROM ),
      .O (\bridge/pci_target_unit/fifos/outNextGreyCount [0])
    );
    X_FF \bridge/pci_target_unit/fifos/outGreyCount_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/pci_target_unit/fifos/outGreyCount [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_outTransactionCount<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_outTransactionCount_reg<1> (
      .I (\bridge/pci_target_unit/fifos/outNextGreyCount [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/FFX/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_outTransactionCount<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17685.INIT = 16'hD555;
    X_LUT4 C17685(
      .ADR0 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wclock_nempty_detect85 ),
      .ADR1 (syn19420),
      .ADR2 (syn182538),
      .ADR3 (syn19407),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_empty )
    );
    defparam C19297.INIT = 16'hEFFF;
    X_LUT4 C19297(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR1 (syn19420),
      .ADR2 (syn19407),
      .ADR3 (N12616),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty/FROM ),
      .O (\bridge/pci_target_unit/fifos/portA_enable )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty_reg (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/reg_empty ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR_74 (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17932.INIT = 16'h33CC;
    X_LUT4 C17932(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [2]),
      .O (\bridge/pci_target_unit/fifos/outNextGreyCount [1])
    );
    X_INV \bridge/pci_target_unit/fifos/outGreyCount<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/outGreyCount[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/outGreyCount_reg<1> (
      .I (\bridge/pci_target_unit/fifos/outNextGreyCount [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/out_count_en ),
      .SET (\bridge/pci_target_unit/fifos/outGreyCount[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/outGreyCount [1])
    );
    X_OR2 \bridge/pci_target_unit/fifos/outGreyCount<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/outGreyCount[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/outGreyCount[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17930.INIT = 16'h0FF0;
    X_LUT4 C17930(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [2]),
      .O (\bridge/pci_target_unit/fifos/outNextGreyCount [2])
    );
    X_INV \bridge/pci_target_unit/fifos/outGreyCount<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/outGreyCount[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/outGreyCount_reg<2> (
      .I (\bridge/pci_target_unit/fifos/outNextGreyCount [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/out_count_en ),
      .SET (\bridge/pci_target_unit/fifos/outGreyCount[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/outGreyCount [2])
    );
    X_OR2 \bridge/pci_target_unit/fifos/outGreyCount<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/outGreyCount[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/outGreyCount[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/outGreyCount_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/out_count_en ),
      .SET (\bridge/pci_target_unit/fifos/outGreyCount[3]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/outGreyCount [3])
    );
    X_OR2 \bridge/pci_target_unit/fifos/outGreyCount<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/outGreyCount[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/outGreyCount[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19283.INIT = 16'hCFC0;
    X_LUT4 C19283(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [0]),
      .ADR2 (syn19407),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [0]),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/GROM )
    );
    defparam C19286.INIT = 16'hCFC0;
    X_LUT4 C19286(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [1]),
      .ADR2 (syn19407),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [1]),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_raddr_0<1>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/GROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr [0])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_raddr_0<1>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr [1])
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_raddr_0_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0 [0])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_raddr_0<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_raddr_0_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0 [1])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_raddr_0<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19289.INIT = 16'hE4E4;
    X_LUT4 C19289(
      .ADR0 (syn19407),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [2]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/GROM )
    );
    defparam C19292.INIT = 16'hF0AA;
    X_LUT4 C19292(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [3]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [3]),
      .ADR3 (syn19407),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_raddr_0<3>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/GROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr [2])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_raddr_0<3>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr [3])
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_raddr_0_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0 [2])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_raddr_0<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_raddr_0_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0 [3])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_raddr_0<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19295.INIT = 16'hCCAA;
    X_LUT4 C19295(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [4]),
      .ADR2 (VCC),
      .ADR3 (syn19407),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[4]/GROM )
    );
    defparam C19307.INIT = 16'h0055;
    X_LUT4 C19307(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/empty ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/stretched_empty ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[4]/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_raddr_0<4>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[4]/GROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr [4])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_raddr_0<4>/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[4]/FROM ),
      .O (syn19407)
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_raddr_0_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_raddr_0[4]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_raddr_0[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0 [4])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_raddr_0<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_raddr_0[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19071.INIT = 16'hFFF5;
    X_LUT4 C19071(
      .ADR0 (\CRT/go ),
      .ADR1 (VCC),
      .ADR2 (\CRT/crtc_vblank ),
      .ADR3 (\CRT/crtc_hblank ),
      .O (\CRT/drive_blank_reg160 )
    );
    X_INV \CRT/drive_blank_reg/SRMUX (
      .I (N_RST),
      .O (\CRT/drive_blank_reg/SRNOT )
    );
    X_FF \CRT/drive_blank_reg_reg (
      .I (\CRT/drive_blank_reg160 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/drive_blank_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/drive_blank_reg )
    );
    X_OR2 \CRT/drive_blank_reg/FFY/ASYNC_FF_GSR_OR_75 (
      .I0 (\CRT/drive_blank_reg/SRNOT ),
      .I1 (GSR),
      .O (\CRT/drive_blank_reg/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18079.INIT = 16'hEEAA;
    X_LUT4 C18079(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_control_out [0]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/last_int )
    );
    defparam C19463.INIT = 16'hB800;
    X_LUT4 C19463(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_control_out [0]),
      .ADR1 (syn18908),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/FROM ),
      .O (syn18919)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/last_int ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/FFY/ASYNC_FF_GSR_OR_76 (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17780.INIT = 16'hAA00;
    X_LUT4 C17780(
      .ADR0 (\bridge/pci_target_unit/del_sync/N1235 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn23138),
      .O (\bridge/pci_target_unit/del_sync/C1265/N5 )
    );
    defparam C17781.INIT = 16'hA2AA;
    X_LUT4 C17781(
      .ADR0 (\bridge/pci_target_unit/pcit_if_read_completed_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/same_read_reg ),
      .ADR2 (\bridge/out_bckp_trdy_out ),
      .ADR3 (syn19366),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[0]/FROM )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[0]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/del_sync/comp_cycle_count<0>/XUSED (
      .I (\bridge/pci_target_unit/del_sync/comp_cycle_count[0]/FROM ),
      .O (syn23138)
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<0> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [0])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18110.INIT = 16'hCC00;
    X_LUT4 C18110(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/N140 ),
      .ADR2 (VCC),
      .ADR3 (syn22149),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N5 )
    );
    defparam C18111.INIT = 16'h0010;
    X_LUT4 C18111(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/C707 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending ),
      .ADR3 (syn16935),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/FROM ),
      .O (syn22149)
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<0> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19412.INIT = 16'h0A0A;
    X_LUT4 C19412(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2 ),
      .ADR3 (VCC),
      .O (\bridge/configuration/wb_err_cs_bit10_8[9]/GROM )
    );
    defparam C19384.INIT = 16'hFFF0;
    X_LUT4 C19384(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .O (\bridge/configuration/wb_err_cs_bit10_8[9]/FROM )
    );
    X_INV \bridge/configuration/wb_err_cs_bit10_8<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_cs_bit10_8[9]/SRNOT )
    );
    X_BUF \bridge/configuration/wb_err_cs_bit10_8<9>/YUSED (
      .I (\bridge/configuration/wb_err_cs_bit10_8[9]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_mabort_out )
    );
    X_BUF \bridge/configuration/wb_err_cs_bit10_8<9>/XUSED (
      .I (\bridge/configuration/wb_err_cs_bit10_8[9]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [31])
    );
    X_FF \bridge/configuration/wb_err_cs_bit10_8_reg2<9> (
      .I (\bridge/configuration/wb_err_cs_bit10_8[9]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit10_8[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit10_8 [9])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit10_8<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit10_8[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit10_8[9]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17778.INIT = 16'hCC00;
    X_LUT4 C17778(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/N1237 ),
      .ADR2 (VCC),
      .ADR3 (syn23138),
      .O (\bridge/pci_target_unit/del_sync/C1265/N15 )
    );
    defparam C17777.INIT = 16'hAA00;
    X_LUT4 C17777(
      .ADR0 (\bridge/pci_target_unit/del_sync/N1238 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn23138),
      .O (\bridge/pci_target_unit/del_sync/C1265/N20 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<2> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N15 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [2])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<3> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N20 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [3])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18108.INIT = 16'hA0A0;
    X_LUT4 C18108(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/N142 ),
      .ADR1 (VCC),
      .ADR2 (syn22149),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N15 )
    );
    defparam C18107.INIT = 16'hC0C0;
    X_LUT4 C18107(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/N143 ),
      .ADR2 (syn22149),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N20 )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<2> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N15 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<3> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N20 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18179.INIT = 16'hFFF8;
    X_LUT4 C18179(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/C749 ),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/C707 ),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .ADR3 (syn181426),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C78/N44 )
    );
    defparam C18184.INIT = 16'h1100;
    X_LUT4 C18184(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_control_out [1]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_control_out [0]),
      .ADR2 (VCC),
      .ADR3 (syn16935),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/wishbone_slave/c_state<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/c_state<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/FROM ),
      .O (syn181426)
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/c_state_reg<0> (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/C78/N44 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/c_state<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/c_state[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17776.INIT = 16'hCC00;
    X_LUT4 C17776(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/N1239 ),
      .ADR2 (VCC),
      .ADR3 (syn23138),
      .O (\bridge/pci_target_unit/del_sync/C1265/N25 )
    );
    defparam C17775.INIT = 16'hAA00;
    X_LUT4 C17775(
      .ADR0 (\bridge/pci_target_unit/del_sync/N1240 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn23138),
      .O (\bridge/pci_target_unit/del_sync/C1265/N30 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[5]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<4> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N25 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [4])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<5> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [5])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18106.INIT = 16'h8888;
    X_LUT4 C18106(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/N144 ),
      .ADR1 (syn22149),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N25 )
    );
    defparam C18105.INIT = 16'hC0C0;
    X_LUT4 C18105(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/N145 ),
      .ADR2 (syn22149),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N30 )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<4> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N25 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<5> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [5])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18136.INIT = 16'h3330;
    X_LUT4 C18136(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .ADR3 (syn22076),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C78/N31 )
    );
    defparam C18137.INIT = 16'h0088;
    X_LUT4 C18137(
      .ADR0 (\CRT/ssvga_wbm_if/S_41/cell0 ),
      .ADR1 (syn177324),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [1]),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/wishbone_slave/c_state<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/c_state<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/FROM ),
      .O (syn22076)
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/c_state_reg<1> (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/C78/N31 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/c_state<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/c_state[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18182.INIT = 16'hAA0A;
    X_LUT4 C18182(
      .ADR0 (syn177324),
      .ADR1 (VCC),
      .ADR2 (N12360),
      .ADR3 (syn21870),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C78/N18 )
    );
    defparam C18183.INIT = 16'hFFA0;
    X_LUT4 C18183(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/C707 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/C749 ),
      .ADR3 (syn181426),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/wishbone_slave/c_state<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/c_state<2>/XUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/FROM ),
      .O (syn21870)
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/c_state_reg<2> (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/C78/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/c_state<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/c_state[2]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17774.INIT = 16'hA0A0;
    X_LUT4 C17774(
      .ADR0 (\bridge/pci_target_unit/del_sync/N1241 ),
      .ADR1 (VCC),
      .ADR2 (syn23138),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N35 )
    );
    defparam C17773.INIT = 16'hC0C0;
    X_LUT4 C17773(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/N1242 ),
      .ADR2 (syn23138),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N40 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[7]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<6> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N35 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [6])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<7> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N40 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [7])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18104.INIT = 16'hA0A0;
    X_LUT4 C18104(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/N146 ),
      .ADR1 (VCC),
      .ADR2 (syn22149),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N35 )
    );
    defparam C18103.INIT = 16'hCC00;
    X_LUT4 C18103(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/N147 ),
      .ADR2 (VCC),
      .ADR3 (syn22149),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N40 )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<6> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N35 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [6])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<7> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N40 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [7])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17772.INIT = 16'hAA00;
    X_LUT4 C17772(
      .ADR0 (\bridge/pci_target_unit/del_sync/N1243 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn23138),
      .O (\bridge/pci_target_unit/del_sync/C1265/N45 )
    );
    defparam C17771.INIT = 16'hC0C0;
    X_LUT4 C17771(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/N1244 ),
      .ADR2 (syn23138),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/C1265/N50 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_cycle_count<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[9]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<8> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N45 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [8])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_cycle_count_reg<9> (
      .I (\bridge/pci_target_unit/del_sync/C1265/N50 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count [9])
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_cycle_count<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync/comp_cycle_count[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_cycle_count[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18102.INIT = 16'hA0A0;
    X_LUT4 C18102(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/N148 ),
      .ADR1 (VCC),
      .ADR2 (syn22149),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N45 )
    );
    defparam C18101.INIT = 16'hC0C0;
    X_LUT4 C18101(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/N149 ),
      .ADR2 (syn22149),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/C25/N50 )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<8> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N45 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [8])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_cycle_count_reg<9> (
      .I (\bridge/wishbone_slave_unit/del_sync/C25/N50 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [9])
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18620.INIT = 16'hFFEE;
    X_LUT4 C18620(
      .ADR0 (syn20817),
      .ADR1 (syn180261),
      .ADR2 (VCC),
      .ADR3 (syn20807),
      .O (\bridge/out_bckp_ad_out[10]/GROM )
    );
    defparam C18624.INIT = 16'hA8A0;
    X_LUT4 C18624(
      .ADR0 (syn180250),
      .ADR1 (syn180247),
      .ADR2 (syn180248),
      .ADR3 (syn180240),
      .O (\bridge/out_bckp_ad_out[10]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<10>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[10]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<10>/YUSED (
      .I (\bridge/out_bckp_ad_out[10]/GROM ),
      .O (\bridge/output_backup/C3/N66 )
    );
    X_BUF \bridge/out_bckp_ad_out<10>/XUSED (
      .I (\bridge/out_bckp_ad_out[10]/FROM ),
      .O (syn20807)
    );
    X_FF \bridge/output_backup/ad_out_reg<10> (
      .I (\bridge/out_bckp_ad_out[10]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[10]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [10])
    );
    X_OR2 \bridge/out_bckp_ad_out<10>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[10]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[10]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18610.INIT = 16'hF5A0;
    X_LUT4 C18610(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (VCC),
      .ADR2 (syn20835),
      .ADR3 (syn20841),
      .O (\bridge/out_bckp_ad_out[11]/GROM )
    );
    defparam C18611.INIT = 16'hFCF0;
    X_LUT4 C18611(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [11]),
      .ADR2 (syn180270),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\bridge/out_bckp_ad_out[11]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[11]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<11>/YUSED (
      .I (\bridge/out_bckp_ad_out[11]/GROM ),
      .O (\bridge/output_backup/C3/N72 )
    );
    X_BUF \bridge/out_bckp_ad_out<11>/XUSED (
      .I (\bridge/out_bckp_ad_out[11]/FROM ),
      .O (syn20841)
    );
    X_FF \bridge/output_backup/ad_out_reg<11> (
      .I (\bridge/out_bckp_ad_out[11]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [11])
    );
    X_OR2 \bridge/out_bckp_ad_out<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[11]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18460.INIT = 16'hFFCC;
    X_LUT4 C18460(
      .ADR0 (VCC),
      .ADR1 (syn21197),
      .ADR2 (VCC),
      .ADR3 (syn180720),
      .O (\bridge/out_bckp_ad_out[20]/GROM )
    );
    defparam C18461.INIT = 16'hEEEC;
    X_LUT4 C18461(
      .ADR0 (syn181260),
      .ADR1 (syn180719),
      .ADR2 (syn180707),
      .ADR3 (syn180706),
      .O (\bridge/out_bckp_ad_out[20]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<20>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[20]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<20>/YUSED (
      .I (\bridge/out_bckp_ad_out[20]/GROM ),
      .O (\bridge/output_backup/C3/N126 )
    );
    X_BUF \bridge/out_bckp_ad_out<20>/XUSED (
      .I (\bridge/out_bckp_ad_out[20]/FROM ),
      .O (syn180720)
    );
    X_FF \bridge/output_backup/ad_out_reg<20> (
      .I (\bridge/out_bckp_ad_out[20]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[20]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [20])
    );
    X_OR2 \bridge/out_bckp_ad_out<20>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[20]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[20]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18592.INIT = 16'hFFFE;
    X_LUT4 C18592(
      .ADR0 (syn180336),
      .ADR1 (syn20874),
      .ADR2 (syn20882),
      .ADR3 (syn180337),
      .O (\bridge/out_bckp_ad_out[12]/GROM )
    );
    defparam C18593.INIT = 16'hECCC;
    X_LUT4 C18593(
      .ADR0 (\bridge/conf_latency_tim_out [4]),
      .ADR1 (syn20872),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn17101),
      .O (\bridge/out_bckp_ad_out[12]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<12>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[12]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<12>/YUSED (
      .I (\bridge/out_bckp_ad_out[12]/GROM ),
      .O (\bridge/output_backup/C3/N78 )
    );
    X_BUF \bridge/out_bckp_ad_out<12>/XUSED (
      .I (\bridge/out_bckp_ad_out[12]/FROM ),
      .O (syn180337)
    );
    X_FF \bridge/output_backup/ad_out_reg<12> (
      .I (\bridge/out_bckp_ad_out[12]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[12]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [12])
    );
    X_OR2 \bridge/out_bckp_ad_out<12>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[12]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[12]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18444.INIT = 16'hFFF0;
    X_LUT4 C18444(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn21235),
      .ADR3 (syn180766),
      .O (\bridge/out_bckp_ad_out[21]/GROM )
    );
    defparam C18445.INIT = 16'hFFA8;
    X_LUT4 C18445(
      .ADR0 (syn181260),
      .ADR1 (syn180753),
      .ADR2 (syn180752),
      .ADR3 (syn180765),
      .O (\bridge/out_bckp_ad_out[21]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[21]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<21>/YUSED (
      .I (\bridge/out_bckp_ad_out[21]/GROM ),
      .O (\bridge/output_backup/C3/N132 )
    );
    X_BUF \bridge/out_bckp_ad_out<21>/XUSED (
      .I (\bridge/out_bckp_ad_out[21]/FROM ),
      .O (syn180766)
    );
    X_FF \bridge/output_backup/ad_out_reg<21> (
      .I (\bridge/out_bckp_ad_out[21]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [21])
    );
    X_OR2 \bridge/out_bckp_ad_out<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[21]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18574.INIT = 16'hFFFE;
    X_LUT4 C18574(
      .ADR0 (syn180387),
      .ADR1 (syn20922),
      .ADR2 (syn20913),
      .ADR3 (syn180388),
      .O (\bridge/out_bckp_ad_out[13]/GROM )
    );
    defparam C18575.INIT = 16'hFEFA;
    X_LUT4 C18575(
      .ADR0 (syn20909),
      .ADR1 (syn17120),
      .ADR2 (syn180385),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\bridge/out_bckp_ad_out[13]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[13]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<13>/YUSED (
      .I (\bridge/out_bckp_ad_out[13]/GROM ),
      .O (\bridge/output_backup/C3/N84 )
    );
    X_BUF \bridge/out_bckp_ad_out<13>/XUSED (
      .I (\bridge/out_bckp_ad_out[13]/FROM ),
      .O (syn180388)
    );
    X_FF \bridge/output_backup/ad_out_reg<13> (
      .I (\bridge/out_bckp_ad_out[13]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [13])
    );
    X_OR2 \bridge/out_bckp_ad_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18290.INIT = 16'hFFAA;
    X_LUT4 C18290(
      .ADR0 (syn21601),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn181220),
      .O (\bridge/out_bckp_ad_out[30]/GROM )
    );
    defparam C18291.INIT = 16'hFFF8;
    X_LUT4 C18291(
      .ADR0 (syn181260),
      .ADR1 (syn21585),
      .ADR2 (syn181218),
      .ADR3 (syn181217),
      .O (\bridge/out_bckp_ad_out[30]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<30>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[30]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<30>/YUSED (
      .I (\bridge/out_bckp_ad_out[30]/GROM ),
      .O (\bridge/output_backup/C3/N186 )
    );
    X_BUF \bridge/out_bckp_ad_out<30>/XUSED (
      .I (\bridge/out_bckp_ad_out[30]/FROM ),
      .O (syn181220)
    );
    X_FF \bridge/output_backup/ad_out_reg<30> (
      .I (\bridge/out_bckp_ad_out[30]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[30]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [30])
    );
    X_OR2 \bridge/out_bckp_ad_out<30>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[30]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[30]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18429.INIT = 16'hFFEA;
    X_LUT4 C18429(
      .ADR0 (syn180811),
      .ADR1 (syn181260),
      .ADR2 (syn21259),
      .ADR3 (syn21274),
      .O (\bridge/out_bckp_ad_out[22]/GROM )
    );
    defparam C18433.INIT = 16'h00EA;
    X_LUT4 C18433(
      .ADR0 (syn180806),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [22]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\bridge/out_bckp_ad_out[22]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<22>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[22]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<22>/YUSED (
      .I (\bridge/out_bckp_ad_out[22]/GROM ),
      .O (\bridge/output_backup/C3/N138 )
    );
    X_BUF \bridge/out_bckp_ad_out<22>/XUSED (
      .I (\bridge/out_bckp_ad_out[22]/FROM ),
      .O (syn21274)
    );
    X_FF \bridge/output_backup/ad_out_reg<22> (
      .I (\bridge/out_bckp_ad_out[22]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[22]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [22])
    );
    X_OR2 \bridge/out_bckp_ad_out<22>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[22]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[22]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18556.INIT = 16'hFFCC;
    X_LUT4 C18556(
      .ADR0 (VCC),
      .ADR1 (syn20963),
      .ADR2 (VCC),
      .ADR3 (syn180442),
      .O (\bridge/out_bckp_ad_out[14]/GROM )
    );
    defparam C18557.INIT = 16'hFFEA;
    X_LUT4 C18557(
      .ADR0 (syn180440),
      .ADR1 (syn181260),
      .ADR2 (syn20947),
      .ADR3 (syn180439),
      .O (\bridge/out_bckp_ad_out[14]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<14>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[14]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<14>/YUSED (
      .I (\bridge/out_bckp_ad_out[14]/GROM ),
      .O (\bridge/output_backup/C3/N90 )
    );
    X_BUF \bridge/out_bckp_ad_out<14>/XUSED (
      .I (\bridge/out_bckp_ad_out[14]/FROM ),
      .O (syn180442)
    );
    X_FF \bridge/output_backup/ad_out_reg<14> (
      .I (\bridge/out_bckp_ad_out[14]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[14]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [14])
    );
    X_OR2 \bridge/out_bckp_ad_out<14>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[14]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[14]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18271.INIT = 16'hFFF0;
    X_LUT4 C18271(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn21641),
      .ADR3 (syn181275),
      .O (\bridge/out_bckp_ad_out[31]/GROM )
    );
    defparam C18272.INIT = 16'hFEFC;
    X_LUT4 C18272(
      .ADR0 (syn21625),
      .ADR1 (syn181272),
      .ADR2 (syn181273),
      .ADR3 (syn181260),
      .O (\bridge/out_bckp_ad_out[31]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[31]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<31>/YUSED (
      .I (\bridge/out_bckp_ad_out[31]/GROM ),
      .O (\bridge/output_backup/C3/N192 )
    );
    X_BUF \bridge/out_bckp_ad_out<31>/XUSED (
      .I (\bridge/out_bckp_ad_out[31]/FROM ),
      .O (syn181275)
    );
    X_FF \bridge/output_backup/ad_out_reg<31> (
      .I (\bridge/out_bckp_ad_out[31]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [31])
    );
    X_OR2 \bridge/out_bckp_ad_out<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[31]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18413.INIT = 16'hEE44;
    X_LUT4 C18413(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn21313),
      .ADR2 (VCC),
      .ADR3 (syn21307),
      .O (\bridge/out_bckp_ad_out[23]/GROM )
    );
    defparam C18416.INIT = 16'hECEC;
    X_LUT4 C18416(
      .ADR0 (syn16916),
      .ADR1 (syn180855),
      .ADR2 (syn21298),
      .ADR3 (VCC),
      .O (\bridge/out_bckp_ad_out[23]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[23]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<23>/YUSED (
      .I (\bridge/out_bckp_ad_out[23]/GROM ),
      .O (\bridge/output_backup/C3/N144 )
    );
    X_BUF \bridge/out_bckp_ad_out<23>/XUSED (
      .I (\bridge/out_bckp_ad_out[23]/FROM ),
      .O (syn21307)
    );
    X_FF \bridge/output_backup/ad_out_reg<23> (
      .I (\bridge/out_bckp_ad_out[23]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [23])
    );
    X_OR2 \bridge/out_bckp_ad_out<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[23]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18539.INIT = 16'hFFCC;
    X_LUT4 C18539(
      .ADR0 (VCC),
      .ADR1 (syn21003),
      .ADR2 (VCC),
      .ADR3 (syn180492),
      .O (\bridge/out_bckp_ad_out[15]/GROM )
    );
    defparam C18540.INIT = 16'hFEFC;
    X_LUT4 C18540(
      .ADR0 (syn181260),
      .ADR1 (syn180490),
      .ADR2 (syn180489),
      .ADR3 (syn20987),
      .O (\bridge/out_bckp_ad_out[15]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[15]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<15>/YUSED (
      .I (\bridge/out_bckp_ad_out[15]/GROM ),
      .O (\bridge/output_backup/C3/N96 )
    );
    X_BUF \bridge/out_bckp_ad_out<15>/XUSED (
      .I (\bridge/out_bckp_ad_out[15]/FROM ),
      .O (syn180492)
    );
    X_FF \bridge/output_backup/ad_out_reg<15> (
      .I (\bridge/out_bckp_ad_out[15]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [15])
    );
    X_OR2 \bridge/out_bckp_ad_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18396.INIT = 16'hFFFE;
    X_LUT4 C18396(
      .ADR0 (syn180906),
      .ADR1 (syn180907),
      .ADR2 (syn21346),
      .ADR3 (syn21354),
      .O (\bridge/out_bckp_ad_out[24]/GROM )
    );
    defparam C18401.INIT = 16'h0E0C;
    X_LUT4 C18401(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (syn180899),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [24]),
      .O (\bridge/out_bckp_ad_out[24]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<24>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[24]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<24>/YUSED (
      .I (\bridge/out_bckp_ad_out[24]/GROM ),
      .O (\bridge/output_backup/C3/N150 )
    );
    X_BUF \bridge/out_bckp_ad_out<24>/XUSED (
      .I (\bridge/out_bckp_ad_out[24]/FROM ),
      .O (syn21354)
    );
    X_FF \bridge/output_backup/ad_out_reg<24> (
      .I (\bridge/out_bckp_ad_out[24]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[24]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [24])
    );
    X_OR2 \bridge/out_bckp_ad_out<24>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[24]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[24]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18523.INIT = 16'hFC0C;
    X_LUT4 C18523(
      .ADR0 (VCC),
      .ADR1 (syn21041),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn21035),
      .O (\bridge/out_bckp_ad_out[16]/GROM )
    );
    defparam C18526.INIT = 16'hFCEC;
    X_LUT4 C18526(
      .ADR0 (syn180528),
      .ADR1 (syn180535),
      .ADR2 (syn16916),
      .ADR3 (syn180529),
      .O (\bridge/out_bckp_ad_out[16]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<16>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[16]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<16>/YUSED (
      .I (\bridge/out_bckp_ad_out[16]/GROM ),
      .O (\bridge/output_backup/C3/N102 )
    );
    X_BUF \bridge/out_bckp_ad_out<16>/XUSED (
      .I (\bridge/out_bckp_ad_out[16]/FROM ),
      .O (syn21035)
    );
    X_FF \bridge/output_backup/ad_out_reg<16> (
      .I (\bridge/out_bckp_ad_out[16]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[16]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [16])
    );
    X_OR2 \bridge/out_bckp_ad_out<16>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[16]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[16]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18379.INIT = 16'hFFFE;
    X_LUT4 C18379(
      .ADR0 (syn180961),
      .ADR1 (syn180960),
      .ADR2 (syn21385),
      .ADR3 (syn21396),
      .O (\bridge/out_bckp_ad_out[25]/GROM )
    );
    defparam C18384.INIT = 16'h0E0C;
    X_LUT4 C18384(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (syn180951),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [25]),
      .O (\bridge/out_bckp_ad_out[25]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[25]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<25>/YUSED (
      .I (\bridge/out_bckp_ad_out[25]/GROM ),
      .O (\bridge/output_backup/C3/N156 )
    );
    X_BUF \bridge/out_bckp_ad_out<25>/XUSED (
      .I (\bridge/out_bckp_ad_out[25]/FROM ),
      .O (syn21396)
    );
    X_FF \bridge/output_backup/ad_out_reg<25> (
      .I (\bridge/out_bckp_ad_out[25]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [25])
    );
    X_OR2 \bridge/out_bckp_ad_out<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[25]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18507.INIT = 16'hFFF0;
    X_LUT4 C18507(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn21080),
      .ADR3 (syn180583),
      .O (\bridge/out_bckp_ad_out[17]/GROM )
    );
    defparam C18508.INIT = 16'hEEEC;
    X_LUT4 C18508(
      .ADR0 (syn181260),
      .ADR1 (syn180582),
      .ADR2 (syn180569),
      .ADR3 (syn180570),
      .O (\bridge/out_bckp_ad_out[17]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[17]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<17>/YUSED (
      .I (\bridge/out_bckp_ad_out[17]/GROM ),
      .O (\bridge/output_backup/C3/N108 )
    );
    X_BUF \bridge/out_bckp_ad_out<17>/XUSED (
      .I (\bridge/out_bckp_ad_out[17]/FROM ),
      .O (syn180583)
    );
    X_FF \bridge/output_backup/ad_out_reg<17> (
      .I (\bridge/out_bckp_ad_out[17]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [17])
    );
    X_OR2 \bridge/out_bckp_ad_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17698.INIT = 16'h6666;
    X_LUT4 C17698(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [1]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [0]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/GROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<0>/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/GROM ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [0])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/waddr_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr [1])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<0>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [0])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<0>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[0]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18362.INIT = 16'hDD88;
    X_LUT4 C18362(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn21430),
      .ADR2 (VCC),
      .ADR3 (syn21436),
      .O (\bridge/out_bckp_ad_out[26]/GROM )
    );
    defparam C18363.INIT = 16'hEECC;
    X_LUT4 C18363(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [26]),
      .ADR1 (syn180971),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\bridge/out_bckp_ad_out[26]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<26>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[26]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<26>/YUSED (
      .I (\bridge/out_bckp_ad_out[26]/GROM ),
      .O (\bridge/output_backup/C3/N162 )
    );
    X_BUF \bridge/out_bckp_ad_out<26>/XUSED (
      .I (\bridge/out_bckp_ad_out[26]/FROM ),
      .O (syn21436)
    );
    X_FF \bridge/output_backup/ad_out_reg<26> (
      .I (\bridge/out_bckp_ad_out[26]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[26]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [26])
    );
    X_OR2 \bridge/out_bckp_ad_out<26>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[26]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[26]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18492.INIT = 16'hFFEC;
    X_LUT4 C18492(
      .ADR0 (syn21104),
      .ADR1 (syn180628),
      .ADR2 (syn181260),
      .ADR3 (syn21119),
      .O (\bridge/out_bckp_ad_out[18]/GROM )
    );
    defparam C18496.INIT = 16'h00F8;
    X_LUT4 C18496(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [18]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn180623),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\bridge/out_bckp_ad_out[18]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<18>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[18]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<18>/YUSED (
      .I (\bridge/out_bckp_ad_out[18]/GROM ),
      .O (\bridge/output_backup/C3/N114 )
    );
    X_BUF \bridge/out_bckp_ad_out<18>/XUSED (
      .I (\bridge/out_bckp_ad_out[18]/FROM ),
      .O (syn21119)
    );
    X_FF \bridge/output_backup/ad_out_reg<18> (
      .I (\bridge/out_bckp_ad_out[18]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[18]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [18])
    );
    X_OR2 \bridge/out_bckp_ad_out<18>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[18]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[18]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_trdy_critical/C52 .INIT = 16'h01FF;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_trdy_critical/C52 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/trdy_w ),
      .ADR2 (N_IRDY),
      .ADR3 
      (\bridge/pci_target_unit/pci_target_sm/pci_target_trdy_critical/syn71 ),
      .O (\bridge/out_bckp_trdy_out/GROM )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_trdy_critical/C53 .INIT = 16'hCCFE;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_trdy_critical/C53 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/trdy_w ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm ),
      .ADR3 (N_FRAME),
      .O (\bridge/out_bckp_trdy_out/FROM )
    );
    X_INV \bridge/out_bckp_trdy_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_trdy_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_trdy_out/YUSED (
      .I (\bridge/out_bckp_trdy_out/GROM ),
      .O (N12472)
    );
    X_BUF \bridge/out_bckp_trdy_out/XUSED (
      .I (\bridge/out_bckp_trdy_out/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/pci_target_trdy_critical/syn71 )
    );
    X_FF \bridge/output_backup/trdy_out_reg (
      .I (\bridge/out_bckp_trdy_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\bridge/out_bckp_trdy_out/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_trdy_out )
    );
    X_OR2 \bridge/out_bckp_trdy_out/FFY/ASYNC_FF_GSR_OR_77 (
      .I0 (\bridge/out_bckp_trdy_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_trdy_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17696.INIT = 16'h3CF0;
    X_LUT4 C17696(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [0]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [1]),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N318 )
    );
    defparam C17695.INIT = 16'h6CCC;
    X_LUT4 C17695(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [0]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [1]),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N319 )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/waddr_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N318 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr [2])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_waddr<3>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFY/RST )
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbr_waddr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/waddr_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N319 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFX/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr [3])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_waddr<3>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFX/RST )
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbr_waddr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFX/RST ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18343.INIT = 16'hFFEC;
    X_LUT4 C18343(
      .ADR0 (syn181260),
      .ADR1 (syn181062),
      .ADR2 (syn21462),
      .ADR3 (syn21479),
      .O (\bridge/out_bckp_ad_out[27]/GROM )
    );
    defparam C18582.INIT = 16'hEE00;
    X_LUT4 C18582(
      .ADR0 (syn180374),
      .ADR1 (syn180373),
      .ADR2 (VCC),
      .ADR3 (syn181260),
      .O (\bridge/out_bckp_ad_out[27]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[27]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<27>/YUSED (
      .I (\bridge/out_bckp_ad_out[27]/GROM ),
      .O (\bridge/output_backup/C3/N168 )
    );
    X_BUF \bridge/out_bckp_ad_out<27>/XUSED (
      .I (\bridge/out_bckp_ad_out[27]/FROM ),
      .O (syn20913)
    );
    X_FF \bridge/output_backup/ad_out_reg<27> (
      .I (\bridge/out_bckp_ad_out[27]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [27])
    );
    X_OR2 \bridge/out_bckp_ad_out<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[27]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18476.INIT = 16'hFA0A;
    X_LUT4 C18476(
      .ADR0 (syn21158),
      .ADR1 (VCC),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn21152),
      .O (\bridge/out_bckp_ad_out[19]/GROM )
    );
    defparam C18479.INIT = 16'hEECC;
    X_LUT4 C18479(
      .ADR0 (syn21143),
      .ADR1 (syn180672),
      .ADR2 (VCC),
      .ADR3 (syn16916),
      .O (\bridge/out_bckp_ad_out[19]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[19]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<19>/YUSED (
      .I (\bridge/out_bckp_ad_out[19]/GROM ),
      .O (\bridge/output_backup/C3/N120 )
    );
    X_BUF \bridge/out_bckp_ad_out<19>/XUSED (
      .I (\bridge/out_bckp_ad_out[19]/FROM ),
      .O (syn21152)
    );
    X_FF \bridge/output_backup/ad_out_reg<19> (
      .I (\bridge/out_bckp_ad_out[19]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [19])
    );
    X_OR2 \bridge/out_bckp_ad_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_ad_enable_critical/C34 .INIT = 16'hCCCE;
    X_LUT4
     \bridge/pci_target_unit/pci_target_sm/pci_target_ad_enable_critical/C34 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/ad_en_w ),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR3 (N_FRAME),
      .O (\bridge/out_bckp_tar_ad_en_out/GROM )
    );
    defparam \bridge/pci_io_mux/ad_en_high_gen/C24 .INIT = 16'h000F;
    X_LUT4 \bridge/pci_io_mux/ad_en_high_gen/C24 (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_mux_tar_ad_en_in ),
      .ADR3 (\bridge/pci_mux_mas_ad_en_in ),
      .O (\bridge/out_bckp_tar_ad_en_out/FROM )
    );
    X_INV \bridge/out_bckp_tar_ad_en_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_tar_ad_en_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_tar_ad_en_out/YUSED (
      .I (\bridge/out_bckp_tar_ad_en_out/GROM ),
      .O (\bridge/pci_mux_tar_ad_en_in )
    );
    X_BUF \bridge/out_bckp_tar_ad_en_out/XUSED (
      .I (\bridge/out_bckp_tar_ad_en_out/FROM ),
      .O (N12338)
    );
    X_FF \bridge/output_backup/tar_ad_en_out_reg (
      .I (\bridge/out_bckp_tar_ad_en_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/out_bckp_tar_ad_en_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_tar_ad_en_out )
    );
    X_OR2 \bridge/out_bckp_tar_ad_en_out/FFY/ASYNC_FF_GSR_OR_78 (
      .I0 (\bridge/out_bckp_tar_ad_en_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_tar_ad_en_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18325.INIT = 16'hFFFE;
    X_LUT4 C18325(
      .ADR0 (syn181113),
      .ADR1 (syn181114),
      .ADR2 (syn21511),
      .ADR3 (syn21520),
      .O (\bridge/out_bckp_ad_out[28]/GROM )
    );
    defparam C18331.INIT = 16'h3320;
    X_LUT4 C18331(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [28]),
      .ADR3 (syn181107),
      .O (\bridge/out_bckp_ad_out[28]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<28>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[28]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<28>/YUSED (
      .I (\bridge/out_bckp_ad_out[28]/GROM ),
      .O (\bridge/output_backup/C3/N174 )
    );
    X_BUF \bridge/out_bckp_ad_out<28>/XUSED (
      .I (\bridge/out_bckp_ad_out[28]/FROM ),
      .O (syn21520)
    );
    X_FF \bridge/output_backup/ad_out_reg<28> (
      .I (\bridge/out_bckp_ad_out[28]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[28]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [28])
    );
    X_OR2 \bridge/out_bckp_ad_out<28>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[28]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[28]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17693.INIT = 16'h33CC;
    X_LUT4 C17693(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [4]),
      .ADR2 (VCC),
      .ADR3 (syn23454),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N320 )
    );
    defparam C17694.INIT = 16'h8000;
    X_LUT4 C17694(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [0]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [3]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [1]),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_waddr<4>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FROM ),
      .O (syn23454)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/waddr_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N320 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr [4])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_waddr<4>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FFY/RST )
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbr_waddr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[4]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18308.INIT = 16'hFFFE;
    X_LUT4 C18308(
      .ADR0 (syn181166),
      .ADR1 (syn181165),
      .ADR2 (syn21552),
      .ADR3 (syn21560),
      .O (\bridge/out_bckp_ad_out[29]/GROM )
    );
    defparam C18313.INIT = 16'h00F8;
    X_LUT4 C18313(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [29]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn181158),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\bridge/out_bckp_ad_out[29]/FROM )
    );
    X_INV \bridge/out_bckp_ad_out<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_ad_out[29]/SRNOT )
    );
    X_BUF \bridge/out_bckp_ad_out<29>/YUSED (
      .I (\bridge/out_bckp_ad_out[29]/GROM ),
      .O (\bridge/output_backup/C3/N180 )
    );
    X_BUF \bridge/out_bckp_ad_out<29>/XUSED (
      .I (\bridge/out_bckp_ad_out[29]/FROM ),
      .O (syn21560)
    );
    X_FF \bridge/output_backup/ad_out_reg<29> (
      .I (\bridge/out_bckp_ad_out[29]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/output_backup/data_load ),
      .SET (GND),
      .RST (\bridge/out_bckp_ad_out[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_ad_out [29])
    );
    X_OR2 \bridge/out_bckp_ad_out<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/out_bckp_ad_out[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_ad_out[29]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17692.INIT = 16'h6C6C;
    X_LUT4 C17692(
      .ADR0 (syn23454),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [5]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [4]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N321 )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/waddr_reg<5> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N321 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbr_waddr[5]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr [5])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_waddr<5>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[5]/FFY/RST )
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbr_waddr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr[5]/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18143.INIT = 16'h8000;
    X_LUT4 C18143(
      .ADR0 (syn181522),
      .ADR1 (syn181521),
      .ADR2 (syn181520),
      .ADR3 (syn181523),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/wdel_addr_hit )
    );
    defparam C18144.INIT = 16'h8000;
    X_LUT4 C18144(
      .ADR0 (syn181508),
      .ADR1 (syn181511),
      .ADR2 (syn181509),
      .ADR3 (syn181510),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/XUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/FROM ),
      .O (syn181523)
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit_reg (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/wdel_addr_hit ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit )
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/FFY/ASYNC_FF_GSR_OR_79 (
      .I0 (\bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18024.INIT = 16'hC0C0;
    X_LUT4 C18024(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [0]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C25/N6 )
    );
    defparam C18023.INIT = 16'hA0A0;
    X_LUT4 C18023(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [1]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C25/N12 )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[1]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_byte_address_reg<0> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C25/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12594),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_byte_address_reg<1> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C25/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (N12594),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18071.INIT = 16'hFAF8;
    X_LUT4 C18071(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR1 (syn18863),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (syn181624),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C20/N6 )
    );
    defparam C19397.INIT = 16'hA0A8;
    X_LUT4 C19397(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR1 (syn178711),
      .ADR2 (syn178714),
      .ADR3 (syn18863),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/FROM ),
      .O (syn19085)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C20/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/FFY/ASYNC_FF_GSR_OR_80 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req/FFY/ASYNC_FF_GSR_OR )

    );
    defparam \bridge/parity_checker/perr_crit_gen/C40 .INIT = 16'h99FF;
    X_LUT4 \bridge/parity_checker/perr_crit_gen/C40 (
      .ADR0 (N_PAR),
      .ADR1 (\bridge/parity_checker/non_critical_par ),
      .ADR2 (VCC),
      .ADR3 (\bridge/parity_checker/perr_generate ),
      .O (\bridge/out_bckp_perr_out/GROM )
    );
    defparam \bridge/parity_checker/C1138 .INIT = 16'h0002;
    X_LUT4 \bridge/parity_checker/C1138 (
      .ADR0 (\bridge/parity_checker/syn415 ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (\bridge/output_backup/mas_ad_en_out ),
      .ADR3 (\bridge/out_bckp_par_en_out ),
      .O (\bridge/out_bckp_perr_out/FROM )
    );
    X_INV \bridge/out_bckp_perr_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_perr_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_perr_out/YUSED (
      .I (\bridge/out_bckp_perr_out/GROM ),
      .O (N12031)
    );
    X_BUF \bridge/out_bckp_perr_out/XUSED (
      .I (\bridge/out_bckp_perr_out/FROM ),
      .O (\bridge/parity_checker/perr_generate )
    );
    X_FF \bridge/output_backup/perr_out_reg (
      .I (\bridge/out_bckp_perr_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\bridge/out_bckp_perr_out/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_perr_out )
    );
    X_OR2 \bridge/out_bckp_perr_out/FFY/ASYNC_FF_GSR_OR_81 (
      .I0 (\bridge/out_bckp_perr_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_perr_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C20034.INIT = 16'h0010;
    X_LUT4 C20034(
      .ADR0 (N12520),
      .ADR1 (N12521),
      .ADR2 (syn177213),
      .ADR3 (N12519),
      .O (\ACK_I/GROM )
    );
    defparam C20033.INIT = 16'hA000;
    X_LUT4 C20033(
      .ADR0 (ADR_O[10]),
      .ADR1 (VCC),
      .ADR2 (N12119),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .O (\ACK_I/FROM )
    );
    X_INV \ACK_I/SRMUX (
      .I (N_RST),
      .O (\ACK_I/SRNOT )
    );
    X_BUF \ACK_I/YUSED (
      .I (\ACK_I/GROM ),
      .O (N12119)
    );
    X_BUF \ACK_I/XUSED (
      .I (\ACK_I/FROM ),
      .O (\CRT/pal_wr_en )
    );
    X_FF \CRT/ssvga_wbs_if/wbs_ack_o_reg (
      .I (\ACK_I/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\ACK_I/FFY/ASYNC_FF_GSR_OR ),
      .O (ACK_I)
    );
    X_OR2 \ACK_I/FFY/ASYNC_FF_GSR_OR_82 (
      .I0 (\ACK_I/SRNOT ),
      .I1 (GSR),
      .O (\ACK_I/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17795.INIT = 16'h22AA;
    X_LUT4 C17795(
      .ADR0 (\bridge/pci_target_unit/del_sync/sync_comp_req_pending ),
      .ADR1 (syn22771),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync_comp_req_pending_out ),
      .O (\bridge/pci_target_unit/del_sync/C4/N5 )
    );
    defparam C17892.INIT = 16'hAA8A;
    X_LUT4 C17892(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (syn19577),
      .ADR2 (\bridge/pci_target_unit/del_sync_comp_req_pending_out ),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_full_out ),
      .O (\bridge/pci_target_unit/del_sync_comp_req_pending_out/FROM )
    );
    X_INV \bridge/pci_target_unit/del_sync_comp_req_pending_out/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_comp_req_pending_out/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/del_sync_comp_req_pending_out/XUSED (
      .I (\bridge/pci_target_unit/del_sync_comp_req_pending_out/FROM ),
      .O (syn16933)
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_req_pending_reg (
      .I (\bridge/pci_target_unit/del_sync/C4/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (N12543),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync_comp_req_pending_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_comp_req_pending_out )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync_comp_req_pending_out/FFY/ASYNC_FF_GSR_OR_83 (
      .I0 (\bridge/pci_target_unit/del_sync_comp_req_pending_out/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync_comp_req_pending_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18128.INIT = 16'hCC44;
    X_LUT4 C18128(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending ),
      .ADR2 (VCC),
      .ADR3 (syn22096),
      .O (\bridge/wishbone_slave_unit/del_sync/C4/N5 )
    );
    defparam C18129.INIT = 16'hFB00;
    X_LUT4 C18129(
      .ADR0 (syn18863),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR2 (syn22093),
      .ADR3 (syn22095),
      .O (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/FROM ),
      .O (syn22096)
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_req_pending_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/C4/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (N12382),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/FFY/ASYNC_FF_GSR_OR_84 (
      .I0 (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17793.INIT = 16'h2233;
    X_LUT4 C17793(
      .ADR0 (\bridge/pci_target_unit/del_sync/req_rty_exp_clr ),
      .ADR1 (\bridge/pci_target_unit/del_sync/req_comp_pending ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/req_rty_exp_reg ),
      .O (N12601)
    );
    X_INV \bridge/pci_target_unit/pcit_if_read_processing_out/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_read_processing_out/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/req_req_pending_reg (
      .I (N12601),
      .CLK (CLK_BUFGPed),
      .CE (N12544),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pcit_if_read_processing_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_read_processing_out )
    );
    X_OR2
     \bridge/pci_target_unit/pcit_if_read_processing_out/FFY/ASYNC_FF_GSR_OR_85 (
      .I0 (\bridge/pci_target_unit/pcit_if_read_processing_out/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pcit_if_read_processing_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18125.INIT = 16'h5151;
    X_LUT4 C18125(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr ),
      .ADR3 (VCC),
      .O (N12591)
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_req_req_pending_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/req_req_pending_reg (
      .I (N12591),
      .CLK (CLK_BUFGPed),
      .CE (N12383),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_req_req_pending_out/FFY/ASYNC_FF_GSR_OR_86 (
      .I0 (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18198.INIT = 16'h3F2A;
    X_LUT4 C18198(
      .ADR0 (syn181403),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_control_out [0]),
      .ADR2 (syn19088),
      .ADR3 (syn181402),
      .O (\bridge/wishbone_slave_unit/fifos/C2/N5 )
    );
    X_INV \bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_transaction_ready_out_reg (
      .I (\bridge/wishbone_slave_unit/fifos/C2/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out/FFY/ASYNC_FF_GSR_OR_87 (
      .I0 (\bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17914.INIT = 16'hB0F4;
    X_LUT4 C17914(
      .ADR0 (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .ADR1 (\bridge/pci_target_unit/del_sync/req_comp_pending ),
      .ADR2 (\bridge/pci_target_unit/pcit_if_norm_access_to_config_out ),
      .ADR3 (syn19075),
      .O (\bridge/pci_target_unit/pci_target_sm/read_progress )
    );
    defparam C19407.INIT = 16'h0505;
    X_LUT4 C19407(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/pci_target_sm/rd_progress/FROM )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/rd_progress/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/rd_progress/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/rd_progress/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/rd_progress/FROM ),
      .O (syn19075)
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/rd_progress_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/read_progress ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/rd_progress/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/rd_progress )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/rd_progress/FFY/ASYNC_FF_GSR_OR_88 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/rd_progress/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/rd_progress/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19321.INIT = 16'h8800;
    X_LUT4 C19321(
      .ADR0 (syn178849),
      .ADR1 (syn178848),
      .ADR2 (VCC),
      .ADR3 (syn178853),
      .O (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/GROM )
    );
    defparam C19322.INIT = 16'h9000;
    X_LUT4 C19322(
      .ADR0 (\bridge/conf_pci_ba0_out [12]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .ADR2 (syn178847),
      .ADR3 (syn178850),
      .O (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/FROM )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_norm_access_to_config_out )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/FROM ),
      .O (syn178853)
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/FFY/ASYNC_FF_GSR_OR_89 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C18250.INIT = 16'h55AA;
    X_LUT4 C18250(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr [1]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [0]),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [0])
    );
    defparam C18249.INIT = 16'h6666;
    X_LUT4 C18249(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr [1]),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [1])
    );
    X_INV \CRT/ssvga_fifo/sync_gray_rd_ptr<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[1]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<0> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [0]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [0])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<1> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [1]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [1])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18248.INIT = 16'h0FF0;
    X_LUT4 C18248(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [2]),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [3]),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [2])
    );
    defparam C18247.INIT = 16'h0FF0;
    X_LUT4 C18247(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [3]),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [4]),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [3])
    );
    X_INV \CRT/ssvga_fifo/sync_gray_rd_ptr<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[3]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<2> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [2]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [2])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<3> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [3]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [3])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18246.INIT = 16'h5A5A;
    X_LUT4 C18246(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr [5]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [4]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [4])
    );
    defparam C18245.INIT = 16'h3C3C;
    X_LUT4 C18245(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr [5]),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [6]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [5])
    );
    X_INV \CRT/ssvga_fifo/sync_gray_rd_ptr<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[5]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<4> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [4]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [4])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<5> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [5]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [5])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18244.INIT = 16'h55AA;
    X_LUT4 C18244(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [6]),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [6])
    );
    defparam C18243.INIT = 16'h55AA;
    X_LUT4 C18243(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [8]),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [7])
    );
    X_INV \CRT/ssvga_fifo/sync_gray_rd_ptr<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[7]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<6> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [6]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [6])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<7> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [7]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [7])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/C1120 .INIT = 16'h3300;
    X_LUT4 \bridge/parity_checker/C1120 (
      .ADR0 (VCC),
      .ADR1 (\bridge/out_bckp_frame_en_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/in_reg_frame_out ),
      .O (\bridge/parity_checker/frame_dec2201 )
    );
    defparam C19218.INIT = 16'h3030;
    X_LUT4 C19218(
      .ADR0 (VCC),
      .ADR1 (\bridge/in_reg_frame_out ),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/FROM )
    );
    X_INV \bridge/pci_target_unit/del_sync/req_rty_exp_clr/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/del_sync/req_rty_exp_clr/XUSED (
      .I (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_control_out[2] )
    );
    X_FF \bridge/parity_checker/frame_dec2_reg (
      .I (\bridge/parity_checker/frame_dec2201 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/parity_checker/frame_dec2 )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/req_rty_exp_clr/FFY/ASYNC_FF_GSR_OR_90 (
      .I0 (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/req_rty_exp_clr_reg (
      .I (\bridge/pci_target_unit/del_sync/req_rty_exp_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_clr )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/req_rty_exp_clr/FFX/ASYNC_FF_GSR_OR_91 (
      .I0 (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_clr/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18242.INIT = 16'h3C3C;
    X_LUT4 C18242(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr [8]),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [9]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/gray_rd_ptr [8])
    );
    defparam C20007.INIT = 16'hBB88;
    X_LUT4 C20007(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr_plus1 [8]),
      .ADR1 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [8]),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FROM )
    );
    X_INV \CRT/ssvga_fifo/sync_gray_rd_ptr<9>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/SRNOT )
    );
    X_BUF \CRT/ssvga_fifo/sync_gray_rd_ptr<9>/XUSED (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FROM ),
      .O (\CRT/ssvga_fifo/C6/N48 )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<8> (
      .I (\CRT/ssvga_fifo/gray_rd_ptr [8]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [8])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/read_ptr_sync/sync_data_out_reg<9> (
      .I (\CRT/ssvga_fifo/rd_ptr [9]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr [9])
    );
    X_OR2 \CRT/ssvga_fifo/sync_gray_rd_ptr<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/sync_gray_rd_ptr[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17715.INIT = 16'h6666;
    X_LUT4 C17715(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [1]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [1])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [1])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<1>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[1]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[1]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17703.INIT = 16'h6666;
    X_LUT4 C17703(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [3]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [2])
    );
    defparam C17712.INIT = 16'h55AA;
    X_LUT4 C17712(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [4]),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [3])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [2])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<3>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [3])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<3>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17699.INIT = 16'h0FF0;
    X_LUT4 C17699(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [4]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [5]),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [4])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/calc_wgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [4])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<5>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next_reg<5> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_waddr [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [5])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<5>/FFX/SETOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFX/SET )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFX/SET ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next[5]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17896.INIT = 16'hEEEE;
    X_LUT4 C17896(
      .ADR0 (ACK_I),
      .ADR1 (ERR_I),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt379 )
    );
    defparam C18820.INIT = 16'h00CC;
    X_LUT4 C18820(
      .ADR0 (VCC),
      .ADR1 (ERR_I),
      .ADR2 (VCC),
      .ADR3 (ACK_I),
      .O (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt/FROM )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/reset_rty_cnt/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/reset_rty_cnt/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C1183 )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/reset_rty_cnt_reg (
      .I (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt379 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt )
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/reset_rty_cnt/FFY/ASYNC_FF_GSR_OR_92 (
      .I0 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18004.INIT = 16'hFF80;
    X_LUT4 C18004(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [10]),
      .ADR2 (N12594),
      .ADR3 (syn181845),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N54 )
    );
    defparam C18005.INIT = 16'h2F20;
    X_LUT4 C18005(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [10]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3392 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[10]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<10>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[10]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<10>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[10]/FROM ),
      .O (syn181845)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<10> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N54 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[10]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [10])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<10>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[10]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[10]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18002.INIT = 16'hFF80;
    X_LUT4 C18002(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [11]),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (syn181850),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N60 )
    );
    defparam C18003.INIT = 16'h4F40;
    X_LUT4 C18003(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [11]),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3393 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[11]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[11]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<11>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[11]/FROM ),
      .O (syn181850)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<11> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N60 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [11])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[11]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17984.INIT = 16'hFF80;
    X_LUT4 C17984(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [20]),
      .ADR3 (syn181895),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N114 )
    );
    defparam C17985.INIT = 16'h0CAC;
    X_LUT4 C17985(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [20]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3402 ),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[20]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<20>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[20]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<20>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[20]/FROM ),
      .O (syn181895)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<20> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N114 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[20]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [20])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<20>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[20]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[20]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18000.INIT = 16'hFF80;
    X_LUT4 C18000(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [12]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (syn181855),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N66 )
    );
    defparam C18001.INIT = 16'h0ACA;
    X_LUT4 C18001(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3394 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [12]),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[12]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<12>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[12]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<12>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[12]/FROM ),
      .O (syn181855)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<12> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N66 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[12]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [12])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<12>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[12]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[12]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/serr_crit_gen/C32 .INIT = 16'hF9FF;
    X_LUT4 \bridge/parity_checker/serr_crit_gen/C32 (
      .ADR0 (N_PAR),
      .ADR1 (\bridge/parity_checker/non_critical_par ),
      .ADR2 (\bridge/in_reg_frame_out ),
      .ADR3 (\bridge/parity_checker/frame_dec2 ),
      .O (\bridge/parity_checker/pci_perr_en_reg/GROM )
    );
    defparam \bridge/parity_checker/perr_en_crit_gen/C72 .INIT = 16'h0880;
    X_LUT4 \bridge/parity_checker/perr_en_crit_gen/C72 (
      .ADR0 (\bridge/conf_perr_response_out ),
      .ADR1 (\bridge/parity_checker/perr_generate ),
      .ADR2 (\bridge/parity_checker/non_critical_par ),
      .ADR3 (N_PAR),
      .O (\bridge/parity_checker/perr_en_crit_gen/perr )
    );
    X_INV \bridge/parity_checker/pci_perr_en_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/parity_checker/pci_perr_en_reg/SRNOT )
    );
    X_BUF \bridge/parity_checker/pci_perr_en_reg/YUSED (
      .I (\bridge/parity_checker/pci_perr_en_reg/GROM ),
      .O (N12029)
    );
    X_FF \bridge/output_backup/serr_out_reg (
      .I (\bridge/parity_checker/pci_perr_en_reg/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\bridge/parity_checker/pci_perr_en_reg/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_serr_out )
    );
    X_OR2 \bridge/parity_checker/pci_perr_en_reg/FFY/ASYNC_FF_GSR_OR_93 (
      .I0 (\bridge/parity_checker/pci_perr_en_reg/SRNOT ),
      .I1 (GSR),
      .O (\bridge/parity_checker/pci_perr_en_reg/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/parity_checker/perr_en_crit_gen/perr_en_reg_out_reg (
      .I (\bridge/parity_checker/perr_en_crit_gen/perr ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/parity_checker/pci_perr_en_reg/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/parity_checker/pci_perr_en_reg )
    );
    X_OR2 \bridge/parity_checker/pci_perr_en_reg/FFX/ASYNC_FF_GSR_OR_94 (
      .I0 (\bridge/parity_checker/pci_perr_en_reg/SRNOT ),
      .I1 (GSR),
      .O (\bridge/parity_checker/pci_perr_en_reg/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17982.INIT = 16'hFF80;
    X_LUT4 C17982(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [21]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (syn181900),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N120 )
    );
    defparam C17983.INIT = 16'h5D08;
    X_LUT4 C17983(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [21]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3403 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[21]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[21]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<21>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[21]/FROM ),
      .O (syn181900)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<21> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N120 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [21])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[21]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17998.INIT = 16'hFF80;
    X_LUT4 C17998(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [13]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (syn181860),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N72 )
    );
    defparam C17999.INIT = 16'h7520;
    X_LUT4 C17999(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [13]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3395 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[13]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[13]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<13>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[13]/FROM ),
      .O (syn181860)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<13> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N72 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [13])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17964.INIT = 16'hFF80;
    X_LUT4 C17964(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [30]),
      .ADR3 (syn181945),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N174 )
    );
    defparam C17965.INIT = 16'h30B8;
    X_LUT4 C17965(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [30]),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3412 ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[30]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<30>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[30]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<30>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[30]/FROM ),
      .O (syn181945)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<30> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N174 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[30]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [30])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<30>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[30]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[30]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17980.INIT = 16'hFF80;
    X_LUT4 C17980(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [22]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (syn181905),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N126 )
    );
    defparam C17981.INIT = 16'h7250;
    X_LUT4 C17981(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3404 ),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [22]),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[22]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<22>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[22]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<22>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[22]/FROM ),
      .O (syn181905)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<22> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N126 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[22]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [22])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<22>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[22]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[22]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17996.INIT = 16'hFF80;
    X_LUT4 C17996(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [14]),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (syn181865),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N78 )
    );
    defparam C17997.INIT = 16'h7520;
    X_LUT4 C17997(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [14]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3396 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[14]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<14>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[14]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<14>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[14]/FROM ),
      .O (syn181865)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<14> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N78 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[14]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [14])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<14>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[14]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[14]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17962.INIT = 16'hFF80;
    X_LUT4 C17962(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [31]),
      .ADR2 (N12594),
      .ADR3 (syn181950),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N180 )
    );
    defparam C17963.INIT = 16'h5C0C;
    X_LUT4 C17963(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3413 ),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [31]),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[31]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[31]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<31>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[31]/FROM ),
      .O (syn181950)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<31> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N180 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [31])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[31]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17978.INIT = 16'hFF80;
    X_LUT4 C17978(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [23]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (syn181910),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N132 )
    );
    defparam C17979.INIT = 16'h4F40;
    X_LUT4 C17979(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [23]),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3405 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[23]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[23]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<23>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[23]/FROM ),
      .O (syn181910)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<23> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N132 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [23])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[23]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17994.INIT = 16'hFF80;
    X_LUT4 C17994(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [15]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (syn181870),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N84 )
    );
    defparam C17995.INIT = 16'h2E22;
    X_LUT4 C17995(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3397 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [15]),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[15]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[15]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<15>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[15]/FROM ),
      .O (syn181870)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<15> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N84 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [15])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17976.INIT = 16'hFF80;
    X_LUT4 C17976(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [24]),
      .ADR3 (syn181915),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N138 )
    );
    defparam C17977.INIT = 16'h22F0;
    X_LUT4 C17977(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [24]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3406 ),
      .ADR3 (N12594),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[24]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<24>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[24]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<24>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[24]/FROM ),
      .O (syn181915)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<24> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N138 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[24]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [24])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<24>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[24]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[24]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17992.INIT = 16'hFF80;
    X_LUT4 C17992(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [16]),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (syn181875),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N90 )
    );
    defparam C17993.INIT = 16'h3B08;
    X_LUT4 C17993(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [16]),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3398 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[16]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<16>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[16]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<16>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[16]/FROM ),
      .O (syn181875)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<16> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N90 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[16]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [16])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<16>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[16]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[16]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17974.INIT = 16'hFF80;
    X_LUT4 C17974(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [25]),
      .ADR3 (syn181920),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N144 )
    );
    defparam C17975.INIT = 16'h0CAA;
    X_LUT4 C17975(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3407 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [25]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (N12594),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[25]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[25]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<25>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[25]/FROM ),
      .O (syn181920)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<25> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N144 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [25])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[25]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17990.INIT = 16'hFF80;
    X_LUT4 C17990(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [17]),
      .ADR2 (N12594),
      .ADR3 (syn181880),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N96 )
    );
    defparam C17991.INIT = 16'h50CC;
    X_LUT4 C17991(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3399 ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [17]),
      .ADR3 (N12594),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[17]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[17]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<17>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[17]/FROM ),
      .O (syn181880)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<17> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N96 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [17])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17972.INIT = 16'hFF80;
    X_LUT4 C17972(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [26]),
      .ADR3 (syn181925),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N150 )
    );
    defparam C17973.INIT = 16'h7430;
    X_LUT4 C17973(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3408 ),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [26]),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[26]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<26>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[26]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<26>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[26]/FROM ),
      .O (syn181925)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<26> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N150 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[26]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [26])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<26>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[26]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[26]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17988.INIT = 16'hFF80;
    X_LUT4 C17988(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [18]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (syn181885),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N102 )
    );
    defparam C17989.INIT = 16'h22F0;
    X_LUT4 C17989(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [18]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3400 ),
      .ADR3 (N12594),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[18]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<18>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[18]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<18>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[18]/FROM ),
      .O (syn181885)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<18> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N102 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[18]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [18])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<18>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[18]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[18]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17970.INIT = 16'hFF80;
    X_LUT4 C17970(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [27]),
      .ADR3 (syn181930),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N156 )
    );
    defparam C17971.INIT = 16'h7520;
    X_LUT4 C17971(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [27]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3409 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[27]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[27]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<27>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[27]/FROM ),
      .O (syn181930)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<27> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N156 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [27])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[27]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17986.INIT = 16'hFF80;
    X_LUT4 C17986(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [19]),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR3 (syn181890),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N108 )
    );
    defparam C17987.INIT = 16'h2F20;
    X_LUT4 C17987(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [19]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/N3401 ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[19]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[19]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<19>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[19]/FROM ),
      .O (syn181890)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<19> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N108 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [19])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18033.INIT = 16'hAFAC;
    X_LUT4 C18033(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3190 ),
      .ADR1 (\bridge/conf_cache_line_size_out [0]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/C188 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N6 )
    );
    defparam C18034.INIT = 16'hEFEF;
    X_LUT4 C18034(
      .ADR0 (\bridge/conf_cache_line_size_out [6]),
      .ADR1 (\bridge/conf_cache_line_size_out [7]),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_bc_out [1]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/read_count<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/read_count<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C188 )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<0> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[0]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17968.INIT = 16'hFF80;
    X_LUT4 C17968(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (N12594),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [28]),
      .ADR3 (syn181935),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N162 )
    );
    defparam C17969.INIT = 16'h44F0;
    X_LUT4 C17969(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [28]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3410 ),
      .ADR3 (N12594),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[28]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<28>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[28]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<28>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[28]/FROM ),
      .O (syn181935)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<28> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N162 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[28]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [28])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<28>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[28]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[28]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17966.INIT = 16'hFF80;
    X_LUT4 C17966(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [29]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (N12594),
      .ADR3 (syn181940),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N168 )
    );
    defparam C17967.INIT = 16'h5C0C;
    X_LUT4 C17967(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3411 ),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [29]),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[29]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_address_out<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[29]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_address_out<29>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out[29]/FROM ),
      .O (syn181940)
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/current_dword_address_reg<29> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3276/N168 ),
      .CLK (CLK_BUFGPed),
      .CE (N12436),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out [29])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_address_out<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_address_out[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_address_out[29]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18031.INIT = 16'hCCFA;
    X_LUT4 C18031(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/C188 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3192 ),
      .ADR2 (\bridge/conf_cache_line_size_out [2]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N18 )
    );
    defparam C18030.INIT = 16'hAAFC;
    X_LUT4 C18030(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3193 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/C188 ),
      .ADR2 (\bridge/conf_cache_line_size_out [3]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N24 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/read_count<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<2> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<3> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N24 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18029.INIT = 16'hBBB8;
    X_LUT4 C18029(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3194 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR2 (\bridge/conf_cache_line_size_out [4]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/C188 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N30 )
    );
    defparam C18028.INIT = 16'hDDD8;
    X_LUT4 C18028(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3195 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/C188 ),
      .ADR3 (\bridge/conf_cache_line_size_out [5]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N36 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/read_count<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<4> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<5> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [5])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[5]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17924.INIT = 16'h7878;
    X_LUT4 C17924(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [2]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/N2000 )
    );
    defparam C17923.INIT = 16'h78F0;
    X_LUT4 C17923(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [1]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [0]),
      .O (\bridge/pci_target_unit/fifos/N2001 )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_outTransactionCount<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_outTransactionCount_reg<2> (
      .I (\bridge/pci_target_unit/fifos/N2000 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_outTransactionCount<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_outTransactionCount_reg<3> (
      .I (\bridge/pci_target_unit/fifos/N2001 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/FFX/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_outTransactionCount<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18083.INIT = 16'hECCC;
    X_LUT4 C18083(
      .ADR0 (syn22096),
      .ADR1 (syn22189),
      .ADR2 (N12426),
      .ADR3 (N12594),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C0/N6 )
    );
    defparam C19471.INIT = 16'h0003;
    X_LUT4 C19471(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/FROM ),
      .O (N12594)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/del_read_req_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C0/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/FFY/ASYNC_FF_GSR_OR_95 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18027.INIT = 16'hC0C0;
    X_LUT4 C18027(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3196 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N42 )
    );
    defparam C18026.INIT = 16'hA0A0;
    X_LUT4 C18026(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3197 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N48 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/read_count<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<6> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N42 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [6])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<7> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N48 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [7])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[7]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18091.INIT = 16'hAA00;
    X_LUT4 C18091(
      .ADR0 (syn181605),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn181606),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C17/N5 )
    );
    defparam C18092.INIT = 16'h0001;
    X_LUT4 C18092(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [7]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [6]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [5]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [8]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_bound/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/read_bound/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/read_bound/FROM ),
      .O (syn181606)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_bound_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C17/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST (GSR),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_bound )
    );
    defparam C18025.INIT = 16'hA0A0;
    X_LUT4 C18025(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/N3198 ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N53 )
    );
    defparam C18032.INIT = 16'hAAFC;
    X_LUT4 C18032(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3191 ),
      .ADR1 (\bridge/conf_cache_line_size_out [1]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/C188 ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N12 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/read_count<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<8> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N53 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [8])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/read_count_reg<1> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C3277/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (N12466),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/read_count<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/read_count[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17756.INIT = 16'h5A5A;
    X_LUT4 C17756(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [1]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next [1])
    );
    defparam \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<1>/F .INIT = 16'h0000;
    X_LUT4 \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<1>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/FROM ),
      .O (GLOBAL_LOGIC0_6)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17735.INIT = 16'h55AA;
    X_LUT4 C17735(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [2]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next [2])
    );
    defparam C17752.INIT = 16'h33CC;
    X_LUT4 C17752(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [3]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [4]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next [3])
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/calc_wgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19037.INIT = 16'hFFD5;
    X_LUT4 C19037(
      .ADR0 (N_LED),
      .ADR1 (\CRT/ssvga_fifo/S_28/cell0 ),
      .ADR2 (\CRT/go ),
      .ADR3 (syn20069),
      .O (\CRT/ssvga_wbm_if/frame_read_in )
    );
    defparam C19038.INIT = 16'h8000;
    X_LUT4 C19038(
      .ADR0 (\CRT/fifo_wr_en ),
      .ADR1 (syn179377),
      .ADR2 (syn179378),
      .ADR3 (syn179382),
      .O (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FROM ),
      .O (syn20069)
    );
    X_FF \CRT/ssvga_wbm_if/frame_read_reg (
      .I (\CRT/ssvga_wbm_if/frame_read_in ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FFY/ASYNC_FF_GSR_OR )
,
      .O (\CRT/ssvga_wbm_if/frame_read )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FFY/ASYNC_FF_GSR_OR_96 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FFX/ASYNC_FF_GSR_OR_97 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17912.INIT = 16'h0001;
    X_LUT4 C17912(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_full_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_two_left_out ),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_full ),
      .O (\bridge/pci_target_unit/pci_target_sm/write_to_fifo )
    );
    defparam C17915.INIT = 16'h3020;
    X_LUT4 C17915(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .ADR2 (\bridge/pci_target_unit/del_sync/req_comp_pending ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty ),
      .O (\bridge/pci_target_unit/pci_target_sm/read_from_fifo )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/rd_from_fifo/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/wr_to_fifo_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/write_to_fifo ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/wr_to_fifo )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/rd_from_fifo/FFY/ASYNC_FF_GSR_OR_98 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/rd_from_fifo_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/read_from_fifo ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/rd_from_fifo/FFX/ASYNC_FF_GSR_OR_99 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18940.INIT = 16'hCC00;
    X_LUT4 C18940(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/N326 ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/cell25 ),
      .O (\CRT/ssvga_crtc/C532/N5 )
    );
    defparam C18941.INIT = 16'hF7FF;
    X_LUT4 C18941(
      .ADR0 (\CRT/ssvga_crtc/vcntr [1]),
      .ADR1 (syn179548),
      .ADR2 (syn179572),
      .ADR3 (\CRT/ssvga_crtc/vcntr [4]),
      .O (\CRT/ssvga_crtc/vcntr[0]/FROM )
    );
    X_INV \CRT/ssvga_crtc/vcntr<0>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/vcntr[0]/SRNOT )
    );
    X_BUF \CRT/ssvga_crtc/vcntr<0>/XUSED (
      .I (\CRT/ssvga_crtc/vcntr[0]/FROM ),
      .O (\CRT/ssvga_crtc/cell25 )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<0> (
      .I (\CRT/ssvga_crtc/C532/N5 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [0])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[0]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18938.INIT = 16'h8888;
    X_LUT4 C18938(
      .ADR0 (\CRT/ssvga_crtc/cell25 ),
      .ADR1 (\CRT/ssvga_crtc/N327 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/C532/N10 )
    );
    X_INV \CRT/ssvga_crtc/vcntr<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/vcntr[1]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<1> (
      .I (\CRT/ssvga_crtc/C532/N10 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [1])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18937.INIT = 16'hAA00;
    X_LUT4 C18937(
      .ADR0 (\CRT/ssvga_crtc/cell25 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/N328 ),
      .O (\CRT/ssvga_crtc/C532/N15 )
    );
    defparam C18936.INIT = 16'hA0A0;
    X_LUT4 C18936(
      .ADR0 (\CRT/ssvga_crtc/cell25 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/N329 ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/C532/N20 )
    );
    X_INV \CRT/ssvga_crtc/vcntr<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/vcntr[3]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<2> (
      .I (\CRT/ssvga_crtc/C532/N15 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [2])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<3> (
      .I (\CRT/ssvga_crtc/C532/N20 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [3])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18935.INIT = 16'hC0C0;
    X_LUT4 C18935(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/cell25 ),
      .ADR2 (\CRT/ssvga_crtc/N330 ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/C532/N25 )
    );
    defparam C18934.INIT = 16'hAA00;
    X_LUT4 C18934(
      .ADR0 (\CRT/ssvga_crtc/cell25 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/N331 ),
      .O (\CRT/ssvga_crtc/C532/N30 )
    );
    X_INV \CRT/ssvga_crtc/vcntr<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/vcntr[5]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<4> (
      .I (\CRT/ssvga_crtc/C532/N25 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [4])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<5> (
      .I (\CRT/ssvga_crtc/C532/N30 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [5])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18933.INIT = 16'hA0A0;
    X_LUT4 C18933(
      .ADR0 (\CRT/ssvga_crtc/N332 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/cell25 ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/C532/N35 )
    );
    defparam C18932.INIT = 16'hC0C0;
    X_LUT4 C18932(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/N333 ),
      .ADR2 (\CRT/ssvga_crtc/cell25 ),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/C532/N40 )
    );
    X_INV \CRT/ssvga_crtc/vcntr<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/vcntr[7]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<6> (
      .I (\CRT/ssvga_crtc/C532/N35 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [6])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<7> (
      .I (\CRT/ssvga_crtc/C532/N40 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [7])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18077.INIT = 16'hFCFC;
    X_LUT4 C18077(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/write_req_int327 )
    );
    defparam C18088.INIT = 16'hCC08;
    X_LUT4 C18088(
      .ADR0 (syn19064),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 ),
      .ADR3 (syn18863),
      .O (syn22180)
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/write_req_int_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/write_req_int327 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/write_req_int )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/FFY/ASYNC_FF_GSR_OR_100 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/del_write_req_reg (
      .I (syn22180),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/FFX/ASYNC_FF_GSR_OR_101 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18931.INIT = 16'hAA00;
    X_LUT4 C18931(
      .ADR0 (\CRT/ssvga_crtc/cell25 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/N334 ),
      .O (\CRT/ssvga_crtc/C532/N45 )
    );
    defparam C18930.INIT = 16'hAA00;
    X_LUT4 C18930(
      .ADR0 (\CRT/ssvga_crtc/cell25 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/N335 ),
      .O (\CRT/ssvga_crtc/C532/N50 )
    );
    X_INV \CRT/ssvga_crtc/vcntr<9>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/vcntr[9]/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<8> (
      .I (\CRT/ssvga_crtc/C532/N45 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [8])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/vcntr_reg<9> (
      .I (\CRT/ssvga_crtc/C532/N50 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12152),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/vcntr[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/vcntr [9])
    );
    X_OR2 \CRT/ssvga_crtc/vcntr<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_crtc/vcntr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/vcntr[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19068.INIT = 16'hCC40;
    X_LUT4 C19068(
      .ADR0 (\CRT/ssvga_fifo/S_28/cell0 ),
      .ADR1 (N_LED),
      .ADR2 (\CRT/go ),
      .ADR3 (syn20013),
      .O (\CRT/C0/N5 )
    );
    defparam C19069.INIT = 16'h8800;
    X_LUT4 C19069(
      .ADR0 (\CRT/crtc_hblank ),
      .ADR1 (\CRT/crtc_vblank ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/S_43/cell0 ),
      .O (\CRT/go/FROM )
    );
    X_INV \CRT/go/SRMUX (
      .I (N_RST),
      .O (\CRT/go/SRNOT )
    );
    X_BUF \CRT/go/XUSED (
      .I (\CRT/go/FROM ),
      .O (syn20013)
    );
    X_FF \CRT/go_reg (
      .I (\CRT/C0/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/go/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/go )
    );
    X_OR2 \CRT/go/FFY/ASYNC_FF_GSR_OR_102 (
      .I0 (\CRT/go/SRNOT ),
      .I1 (GSR),
      .O (\CRT/go/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18800.INIT = 16'hAAF0;
    X_LUT4 C18800(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [0]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [0])
      ,
      .ADR3 (syn18908),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/GROM )
    );
    defparam C19464.INIT = 16'h000F;
    X_LUT4 C19464(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/in_reg_devsel_out ),
      .ADR3 (\bridge/in_reg_trdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<0>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [0])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/FROM ),
      .O (syn18908)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [0])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18759.INIT = 16'hFC30;
    X_LUT4 C18759(
      .ADR0 (VCC),
      .ADR1 (syn18908),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [1])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [1]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[1]/GROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[1]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<1>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[1]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [1])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<1> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [1])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18746.INIT = 16'hF3C0;
    X_LUT4 C18746(
      .ADR0 (VCC),
      .ADR1 (syn18908),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [2]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [2])
      ,
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/GROM )
    );
    defparam C18733.INIT = 16'hFC0C;
    X_LUT4 C18733(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [3])
      ,
      .ADR2 (syn18908),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [3]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<3>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [2])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<3>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [3])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<2> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [2])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<3> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [3])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18714.INIT = 16'hF3C0;
    X_LUT4 C18714(
      .ADR0 (VCC),
      .ADR1 (syn18908),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [4]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [4])
      ,
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/GROM )
    );
    defparam C18700.INIT = 16'hF0CC;
    X_LUT4 C18700(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [5])
      ,
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [5]),
      .ADR3 (syn18908),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<5>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [4])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<5>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [5])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<4> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [4])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<5> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [5])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18994.INIT = 16'hAFAF;
    X_LUT4 C18994(
      .ADR0 (\CRT/ssvga_fifo/N800 ),
      .ADR1 (VCC),
      .ADR2 (N_LED),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C750/N6 )
    );
    defparam C18986.INIT = 16'hCC00;
    X_LUT4 C18986(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/N801 ),
      .ADR2 (VCC),
      .ADR3 (N_LED),
      .O (\CRT/ssvga_fifo/C750/N11 )
    );
    X_INV \CRT/ssvga_fifo/wr_ptr_plus1<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[1]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_plus1_reg<0> (
      .I (\CRT/ssvga_fifo/C750/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (\CRT/ssvga_fifo/wr_ptr_plus1[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1 [0])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr_plus1<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr_plus1[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_plus1_reg<1> (
      .I (\CRT/ssvga_fifo/C750/N11 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr_plus1[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1 [1])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr_plus1<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr_plus1[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_devsel_critical/C52 .INIT = 16'h01FF;
    X_LUT4
     \bridge/pci_target_unit/pci_target_sm/pci_target_devsel_critical/C52 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/devs_w_frm ),
      .ADR1 (N_IRDY),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/devs_w ),
      .ADR3 
      (\bridge/pci_target_unit/pci_target_sm/pci_target_devsel_critical/syn71 ),
      .O (\bridge/out_bckp_devsel_out/GROM )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_devsel_critical/C53 .INIT = 16'hF5F4;
    X_LUT4
     \bridge/pci_target_unit/pci_target_sm/pci_target_devsel_critical/C53 (
      .ADR0 (N_FRAME),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/devs_w_frm ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/devs_w ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy ),
      .O (\bridge/out_bckp_devsel_out/FROM )
    );
    X_INV \bridge/out_bckp_devsel_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_devsel_out/SRNOT )
    );
    X_BUF \bridge/out_bckp_devsel_out/YUSED (
      .I (\bridge/out_bckp_devsel_out/GROM ),
      .O (N12474)
    );
    X_BUF \bridge/out_bckp_devsel_out/XUSED (
      .I (\bridge/out_bckp_devsel_out/FROM ),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/pci_target_devsel_critical/syn71 )
    );
    X_FF \bridge/output_backup/devsel_out_reg (
      .I (\bridge/out_bckp_devsel_out/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\bridge/out_bckp_devsel_out/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/out_bckp_devsel_out )
    );
    X_OR2 \bridge/out_bckp_devsel_out/FFY/ASYNC_FF_GSR_OR_103 (
      .I0 (\bridge/out_bckp_devsel_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_devsel_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18688.INIT = 16'hAFA0;
    X_LUT4 C18688(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [6]),
      .ADR1 (VCC),
      .ADR2 (syn18908),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [6])
      ,
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/GROM )
    );
    defparam C18678.INIT = 16'hFA0A;
    X_LUT4 C18678(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [7])
      ,
      .ADR1 (VCC),
      .ADR2 (syn18908),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [7]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<7>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [6])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<7>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [7])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<6> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [6])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<7> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [7])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18970.INIT = 16'hC0C0;
    X_LUT4 C18970(
      .ADR0 (VCC),
      .ADR1 (N_LED),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [0]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C0/N40 )
    );
    defparam C18969.INIT = 16'h8888;
    X_LUT4 C18969(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr_plus1 [1]),
      .ADR1 (N_LED),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C0/N35 )
    );
    X_INV \CRT/ssvga_fifo/wr_ptr<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/wr_ptr[1]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_reg<0> (
      .I (\CRT/ssvga_fifo/C0/N40 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr [0])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_reg<1> (
      .I (\CRT/ssvga_fifo/C0/N35 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr [1])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18632.INIT = 16'hD8D8;
    X_LUT4 C18632(
      .ADR0 (syn18908),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [10]),
      .ADR2 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [10]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/GROM )
    );
    defparam C18619.INIT = 16'hCFC0;
    X_LUT4 C18619(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [11]),
      .ADR2 (syn18908),
      .ADR3 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [11]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<11>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [10])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<11>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [11])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<10> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [10])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<11> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [11])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18990.INIT = 16'h8888;
    X_LUT4 C18990(
      .ADR0 (\CRT/ssvga_fifo/N802 ),
      .ADR1 (N_LED),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C750/N16 )
    );
    defparam C18989.INIT = 16'hCC00;
    X_LUT4 C18989(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/N803 ),
      .ADR2 (VCC),
      .ADR3 (N_LED),
      .O (\CRT/ssvga_fifo/C750/N21 )
    );
    X_INV \CRT/ssvga_fifo/wr_ptr_plus1<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[3]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_plus1_reg<2> (
      .I (\CRT/ssvga_fifo/C750/N16 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr_plus1[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1 [2])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr_plus1<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr_plus1[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_plus1_reg<3> (
      .I (\CRT/ssvga_fifo/C750/N21 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr_plus1[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1 [3])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr_plus1<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr_plus1[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18668.INIT = 16'hFC30;
    X_LUT4 C18668(
      .ADR0 (VCC),
      .ADR1 (syn18908),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [8])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [8]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/GROM )
    );
    defparam C18648.INIT = 16'hCDC8;
    X_LUT4 C18648(
      .ADR0 (\bridge/in_reg_trdy_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [9])
      ,
      .ADR2 (\bridge/in_reg_devsel_out ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [9]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<9>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [8])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<9>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [9])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<8> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [8])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<9> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [9])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18968.INIT = 16'hF000;
    X_LUT4 C18968(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [2]),
      .ADR3 (N_LED),
      .O (\CRT/ssvga_fifo/C0/N30 )
    );
    defparam C18967.INIT = 16'hC0C0;
    X_LUT4 C18967(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [3]),
      .ADR2 (N_LED),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C0/N25 )
    );
    X_INV \CRT/ssvga_fifo/wr_ptr<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/wr_ptr[3]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_reg<2> (
      .I (\CRT/ssvga_fifo/C0/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr [2])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_reg<3> (
      .I (\CRT/ssvga_fifo/C0/N25 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr [3])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18475.INIT = 16'hFC0C;
    X_LUT4 C18475(
      .ADR0 (VCC),
      .ADR1 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [20]),
      .ADR2 (syn18908),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [20]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/GROM )
    );
    defparam C18459.INIT = 16'hF3C0;
    X_LUT4 C18459(
      .ADR0 (VCC),
      .ADR1 (syn18908),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [21]),
      .ADR3 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [21]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<21>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [20])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<21>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [21])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<20> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [20])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<21> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [21])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[21]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18609.INIT = 16'hCFC0;
    X_LUT4 C18609(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [12]),
      .ADR2 (syn18908),
      .ADR3 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [12]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/GROM )
    );
    defparam C18591.INIT = 16'hFC0C;
    X_LUT4 C18591(
      .ADR0 (VCC),
      .ADR1 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [13]),
      .ADR2 (syn18908),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [13]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<13>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [12])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<13>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [13])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<12> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [12])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<13> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [13])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18992.INIT = 16'hAA00;
    X_LUT4 C18992(
      .ADR0 (\CRT/ssvga_fifo/N804 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (N_LED),
      .O (\CRT/ssvga_fifo/C750/N26 )
    );
    defparam C18987.INIT = 16'h8888;
    X_LUT4 C18987(
      .ADR0 (N_LED),
      .ADR1 (\CRT/ssvga_fifo/N805 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C750/N31 )
    );
    X_INV \CRT/ssvga_fifo/wr_ptr_plus1<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[5]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_plus1_reg<4> (
      .I (\CRT/ssvga_fifo/C750/N26 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr_plus1[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1 [4])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr_plus1<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr_plus1[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_plus1_reg<5> (
      .I (\CRT/ssvga_fifo/C750/N31 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr_plus1[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1 [5])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr_plus1<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr_plus1[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18056.INIT = 16'h3030;
    X_LUT4 C18056(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [10]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N132 )
    );
    defparam C18055.INIT = 16'h3300;
    X_LUT4 C18055(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [11]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N126 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<11>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<10> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N132 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [10])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<11> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N126 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [11])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[11]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18966.INIT = 16'hCC00;
    X_LUT4 C18966(
      .ADR0 (VCC),
      .ADR1 (N_LED),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/wr_ptr_plus1 [4]),
      .O (\CRT/ssvga_fifo/C0/N20 )
    );
    defparam C18965.INIT = 16'hF000;
    X_LUT4 C18965(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [5]),
      .ADR3 (N_LED),
      .O (\CRT/ssvga_fifo/C0/N15 )
    );
    X_INV \CRT/ssvga_fifo/wr_ptr<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/wr_ptr[5]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_reg<4> (
      .I (\CRT/ssvga_fifo/C0/N20 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr [4])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_reg<5> (
      .I (\CRT/ssvga_fifo/C0/N15 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr [5])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18307.INIT = 16'hF0E4;
    X_LUT4 C18307(
      .ADR0 (\bridge/in_reg_devsel_out ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [30]),
      .ADR2 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [30]),
      .ADR3 (\bridge/in_reg_trdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/GROM )
    );
    defparam C18289.INIT = 16'hF0E4;
    X_LUT4 C18289(
      .ADR0 (\bridge/in_reg_devsel_out ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [31]),
      .ADR2 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [31]),
      .ADR3 (\bridge/in_reg_trdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<31>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [30])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<31>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [31])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<30> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [30])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<31> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [31])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[31]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18443.INIT = 16'hF1E0;
    X_LUT4 C18443(
      .ADR0 (\bridge/in_reg_devsel_out ),
      .ADR1 (\bridge/in_reg_trdy_out ),
      .ADR2 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [22]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [22]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/GROM )
    );
    defparam C18428.INIT = 16'hCCD8;
    X_LUT4 C18428(
      .ADR0 (\bridge/in_reg_trdy_out ),
      .ADR1 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [23]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [23]),
      .ADR3 (\bridge/in_reg_devsel_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<23>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [22])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<23>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [23])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<22> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [22])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<23> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [23])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[23]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18573.INIT = 16'hABA8;
    X_LUT4 C18573(
      .ADR0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [14]),
      .ADR1 (\bridge/in_reg_trdy_out ),
      .ADR2 (\bridge/in_reg_devsel_out ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [14]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/GROM )
    );
    defparam C18555.INIT = 16'hF0E2;
    X_LUT4 C18555(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [15]),
      .ADR1 (\bridge/in_reg_trdy_out ),
      .ADR2 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [15]),
      .ADR3 (\bridge/in_reg_devsel_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<15>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [14])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<15>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [15])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<14> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [14])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<15> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [15])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18991.INIT = 16'hA0A0;
    X_LUT4 C18991(
      .ADR0 (\CRT/ssvga_fifo/N806 ),
      .ADR1 (VCC),
      .ADR2 (N_LED),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C750/N36 )
    );
    defparam C18988.INIT = 16'hC0C0;
    X_LUT4 C18988(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/N807 ),
      .ADR2 (N_LED),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C750/N41 )
    );
    X_INV \CRT/ssvga_fifo/wr_ptr_plus1<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[7]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_plus1_reg<6> (
      .I (\CRT/ssvga_fifo/C750/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr_plus1[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1 [6])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr_plus1<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr_plus1[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_plus1_reg<7> (
      .I (\CRT/ssvga_fifo/C750/N41 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr_plus1[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1 [7])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr_plus1<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr_plus1[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18046.INIT = 16'h00AA;
    X_LUT4 C18046(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [20]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N72 )
    );
    defparam C18045.INIT = 16'h4444;
    X_LUT4 C18045(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [21]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N66 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<21>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<20> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N72 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [20])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<21> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N66 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [21])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[21]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18054.INIT = 16'h00F0;
    X_LUT4 C18054(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [12]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N120 )
    );
    defparam C18053.INIT = 16'h00F0;
    X_LUT4 C18053(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [13]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N114 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<13>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<12> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N120 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [12])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<13> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N114 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [13])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[13]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18964.INIT = 16'hCC00;
    X_LUT4 C18964(
      .ADR0 (VCC),
      .ADR1 (N_LED),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/wr_ptr_plus1 [6]),
      .O (\CRT/ssvga_fifo/C0/N10 )
    );
    defparam C18963.INIT = 16'hA0A0;
    X_LUT4 C18963(
      .ADR0 (N_LED),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [7]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C0/N5 )
    );
    X_INV \CRT/ssvga_fifo/wr_ptr<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/wr_ptr[7]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_reg<6> (
      .I (\CRT/ssvga_fifo/C0/N10 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr [6])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/wr_ptr_reg<7> (
      .I (\CRT/ssvga_fifo/C0/N5 ),
      .CLK (CLK_BUFGPed),
      .CE (N12092),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/wr_ptr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/wr_ptr [7])
    );
    X_OR2 \CRT/ssvga_fifo/wr_ptr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/wr_ptr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/wr_ptr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19148.INIT = 16'hCCF0;
    X_LUT4 C19148(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/rd_progress ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/same_read_reg ),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w/GROM )
    );
    defparam C19147.INIT = 16'hEAC0;
    X_LUT4 C19147(
      .ADR0 (syn19914),
      .ADR1 (syn17035),
      .ADR2 (syn19918),
      .ADR3 (syn17012),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/trdy_w/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/trdy_w/GROM ),
      .O (syn19918)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/trdy_w/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/trdy_w/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w )
    );
    defparam C19304.INIT = 16'hFFFB;
    X_LUT4 C19304(
      .ADR0 (syn19385),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/previous_frame ),
      .ADR2 (\bridge/out_bckp_frame_en_out ),
      .ADR3 (\bridge/in_reg_frame_out ),
      .O (\syn17012/GROM )
    );
    defparam C19151.INIT = 16'hC0C0;
    X_LUT4 C19151(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/N59 ),
      .ADR2 (syn24524),
      .ADR3 (VCC),
      .O (\syn17012/FROM )
    );
    X_BUF \syn17012/YUSED (
      .I (\syn17012/GROM ),
      .O (syn24524)
    );
    X_BUF \syn17012/XUSED (
      .I (\syn17012/FROM ),
      .O (syn17012)
    );
    defparam C19317.INIT = 16'h3BCF;
    X_LUT4 C19317(
      .ADR0 (\bridge/in_reg_cbe_out [0]),
      .ADR1 (\bridge/in_reg_cbe_out [3]),
      .ADR2 (\bridge/in_reg_cbe_out [1]),
      .ADR3 (\bridge/in_reg_cbe_out [2]),
      .O (\syn19385/GROM )
    );
    defparam C19316.INIT = 16'hF531;
    X_LUT4 C19316(
      .ADR0 (\bridge/pci_target_unit/pcit_if_norm_access_to_config_out ),
      .ADR1 (syn17031),
      .ADR2 (syn178869),
      .ADR3 (syn19380),
      .O (\syn19385/FROM )
    );
    X_BUF \syn19385/YUSED (
      .I (\syn19385/GROM ),
      .O (syn178869)
    );
    X_BUF \syn19385/XUSED (
      .I (\syn19385/FROM ),
      .O (syn19385)
    );
    defparam C19131.INIT = 16'hAEAA;
    X_LUT4 C19131(
      .ADR0 (syn19968),
      .ADR1 (syn19366),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/same_read_reg ),
      .ADR3 (syn24519),
      .O (\bridge/pci_target_unit/pci_target_sm/stop_w/GROM )
    );
    defparam C19130.INIT = 16'h3100;
    X_LUT4 C19130(
      .ADR0 (syn24524),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR2 (syn179315),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .O (\bridge/pci_target_unit/pci_target_sm/stop_w/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/stop_w/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/stop_w/GROM ),
      .O (syn179315)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/stop_w/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/stop_w/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/stop_w )
    );
    defparam C19159.INIT = 16'h8000;
    X_LUT4 C19159(
      .ADR0 (syn179246),
      .ADR1 (syn179248),
      .ADR2 (syn179247),
      .ADR3 (syn179249),
      .O (\syn17093/GROM )
    );
    defparam C19156.INIT = 16'hFE00;
    X_LUT4 C19156(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/config_access ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_norm_access_to_config_out ),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/decoder1/S_37/cell0 ),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .O (\syn17093/FROM )
    );
    X_BUF \syn17093/YUSED (
      .I (\syn17093/GROM ),
      .O (\bridge/pci_target_unit/pci_target_if/decoder1/S_37/cell0 )
    );
    X_BUF \syn17093/XUSED (
      .I (\syn17093/FROM ),
      .O (syn17093)
    );
    defparam C19161.INIT = 16'h84CC;
    X_LUT4 C19161(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .ADR1 (syn19865),
      .ADR2 (\bridge/conf_pci_ba1_out [18]),
      .ADR3 (\bridge/conf_pci_am1_out [18]),
      .O (\syn179249/GROM )
    );
    defparam C19160.INIT = 16'h9000;
    X_LUT4 C19160(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .ADR1 (\bridge/conf_pci_ba1_out [19]),
      .ADR2 (syn179245),
      .ADR3 (\bridge/conf_pci_am1_out [19]),
      .O (\syn179249/FROM )
    );
    X_BUF \syn179249/YUSED (
      .I (\syn179249/GROM ),
      .O (syn179245)
    );
    X_BUF \syn179249/XUSED (
      .I (\syn179249/FROM ),
      .O (syn179249)
    );
    defparam C19891.INIT = 16'hFFEC;
    X_LUT4 C19891(
      .ADR0 (syn24559),
      .ADR1 (syn17836),
      .ADR2 (\bridge/configuration/status_bit15_11 [15]),
      .ADR3 (syn177532),
      .O (\SDAT_O[31]/GROM )
    );
    defparam C19890.INIT = 16'hFEF0;
    X_LUT4 C19890(
      .ADR0 (syn177519),
      .ADR1 (syn177518),
      .ADR2 (syn177533),
      .ADR3 (syn177524),
      .O (\SDAT_O[31]/FROM )
    );
    X_BUF \SDAT_O<31>/YUSED (
      .I (\SDAT_O[31]/GROM ),
      .O (syn177533)
    );
    X_BUF \SDAT_O<31>/XUSED (
      .I (\SDAT_O[31]/FROM ),
      .O (SDAT_O[31])
    );
    defparam C19939.INIT = 16'hECA0;
    X_LUT4 C19939(
      .ADR0 (\bridge/configuration/pci_err_cs_bit31_24 [31]),
      .ADR1 (\bridge/configuration/pci_tran_addr1 [31]),
      .ADR2 (\bridge/configuration/C2340 ),
      .ADR3 (\bridge/configuration/C2354 ),
      .O (\syn177518/GROM )
    );
    defparam C19938.INIT = 16'hFAFA;
    X_LUT4 C19938(
      .ADR0 (syn177514),
      .ADR1 (VCC),
      .ADR2 (syn177515),
      .ADR3 (VCC),
      .O (\syn177518/FROM )
    );
    X_BUF \syn177518/YUSED (
      .I (\syn177518/GROM ),
      .O (syn177515)
    );
    X_BUF \syn177518/XUSED (
      .I (\syn177518/FROM ),
      .O (syn177518)
    );
    defparam C19947.INIT = 16'hF888;
    X_LUT4 C19947(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/pci_err_addr [31]),
      .ADR2 (\bridge/configuration/C2370 ),
      .ADR3 (\bridge/conf_pci_ba0_out [19]),
      .O (\syn177514/GROM )
    );
    defparam C19946.INIT = 16'hFEFA;
    X_LUT4 C19946(
      .ADR0 (syn17813),
      .ADR1 (\bridge/configuration/wb_err_cs_bit31_24 [31]),
      .ADR2 (syn177511),
      .ADR3 (\bridge/configuration/C2308 ),
      .O (\syn177514/FROM )
    );
    X_BUF \syn177514/YUSED (
      .I (\syn177514/GROM ),
      .O (syn177511)
    );
    X_BUF \syn177514/XUSED (
      .I (\syn177514/FROM ),
      .O (syn177514)
    );
    defparam C19958.INIT = 16'h0800;
    X_LUT4 C19958(
      .ADR0 (syn50321),
      .ADR1 (syn177541),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .O (\bridge/configuration/C2308/GROM )
    );
    defparam C19957.INIT = 16'hC000;
    X_LUT4 C19957(
      .ADR0 (VCC),
      .ADR1 (syn177397),
      .ADR2 (syn177470),
      .ADR3 (syn177396),
      .O (\bridge/configuration/C2308/FROM )
    );
    X_BUF \bridge/configuration/C2308/YUSED (
      .I (\bridge/configuration/C2308/GROM ),
      .O (syn177470)
    );
    X_BUF \bridge/configuration/C2308/XUSED (
      .I (\bridge/configuration/C2308/FROM ),
      .O (\bridge/configuration/C2308 )
    );
    defparam C19973.INIT = 16'h99FF;
    X_LUT4 C19973(
      .ADR0 (\bridge/conf_wb_ba1_out [15]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [27]),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_wb_am1_out [15]),
      .O (\syn177396/GROM )
    );
    defparam C19962.INIT = 16'h8000;
    X_LUT4 C19962(
      .ADR0 (syn60045),
      .ADR1 (syn60044),
      .ADR2 (syn60046),
      .ADR3 (syn60043),
      .O (\syn177396/FROM )
    );
    X_BUF \syn177396/YUSED (
      .I (\syn177396/GROM ),
      .O (syn60046)
    );
    X_BUF \syn177396/XUSED (
      .I (\syn177396/FROM ),
      .O (syn177396)
    );
    defparam C19965.INIT = 16'hC00C;
    X_LUT4 C19965(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_wb_am1_out [19]),
      .ADR2 (\bridge/conf_wb_ba1_out [19]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [31]),
      .O (\syn177397/GROM )
    );
    defparam C19961.INIT = 16'h8000;
    X_LUT4 C19961(
      .ADR0 (syn60047),
      .ADR1 (syn60049),
      .ADR2 (syn177391),
      .ADR3 (syn60048),
      .O (\syn177397/FROM )
    );
    X_BUF \syn177397/YUSED (
      .I (\syn177397/GROM ),
      .O (syn177391)
    );
    X_BUF \syn177397/XUSED (
      .I (\syn177397/FROM ),
      .O (syn177397)
    );
    defparam C19955.INIT = 16'h8000;
    X_LUT4 C19955(
      .ADR0 (syn177563),
      .ADR1 (syn177397),
      .ADR2 (syn50321),
      .ADR3 (syn177396),
      .O (\syn17813/GROM )
    );
    defparam C19953.INIT = 16'h0080;
    X_LUT4 C19953(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [31]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR2 (\bridge/configuration/C3488 ),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .O (\syn17813/FROM )
    );
    X_BUF \syn17813/YUSED (
      .I (\syn17813/GROM ),
      .O (\bridge/configuration/C3488 )
    );
    X_BUF \syn17813/XUSED (
      .I (\syn17813/FROM ),
      .O (syn17813)
    );
    defparam C19951.INIT = 16'h0004;
    X_LUT4 C19951(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR1 (syn84030),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .O (\bridge/configuration/C2370/GROM )
    );
    defparam C19950.INIT = 16'hA000;
    X_LUT4 C19950(
      .ADR0 (syn177397),
      .ADR1 (VCC),
      .ADR2 (syn177403),
      .ADR3 (syn177396),
      .O (\bridge/configuration/C2370/FROM )
    );
    X_BUF \bridge/configuration/C2370/YUSED (
      .I (\bridge/configuration/C2370/GROM ),
      .O (syn177403)
    );
    X_BUF \bridge/configuration/C2370/XUSED (
      .I (\bridge/configuration/C2370/FROM ),
      .O (\bridge/configuration/C2370 )
    );
    defparam C19949.INIT = 16'h0C00;
    X_LUT4 C19949(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .O (\bridge/configuration/C2338/GROM )
    );
    defparam C19948.INIT = 16'h8000;
    X_LUT4 C19948(
      .ADR0 (syn84030),
      .ADR1 (syn177396),
      .ADR2 (syn177475),
      .ADR3 (syn177397),
      .O (\bridge/configuration/C2338/FROM )
    );
    X_BUF \bridge/configuration/C2338/YUSED (
      .I (\bridge/configuration/C2338/GROM ),
      .O (syn177475)
    );
    X_BUF \bridge/configuration/C2338/XUSED (
      .I (\bridge/configuration/C2338/FROM ),
      .O (\bridge/configuration/C2338 )
    );
    defparam C19943.INIT = 16'h0080;
    X_LUT4 C19943(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .O (\bridge/configuration/C2354/GROM )
    );
    defparam C19942.INIT = 16'h1000;
    X_LUT4 C19942(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR2 (syn177485),
      .ADR3 (syn24500),
      .O (\bridge/configuration/C2354/FROM )
    );
    X_BUF \bridge/configuration/C2354/YUSED (
      .I (\bridge/configuration/C2354/GROM ),
      .O (syn177485)
    );
    X_BUF \bridge/configuration/C2354/XUSED (
      .I (\bridge/configuration/C2354/FROM ),
      .O (\bridge/configuration/C2354 )
    );
    defparam C19941.INIT = 16'h0400;
    X_LUT4 C19941(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .O (\bridge/configuration/C2340/GROM )
    );
    defparam C19940.INIT = 16'h0040;
    X_LUT4 C19940(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR1 (syn24500),
      .ADR2 (syn177480),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .O (\bridge/configuration/C2340/FROM )
    );
    X_BUF \bridge/configuration/C2340/YUSED (
      .I (\bridge/configuration/C2340/GROM ),
      .O (syn177480)
    );
    X_BUF \bridge/configuration/C2340/XUSED (
      .I (\bridge/configuration/C2340/FROM ),
      .O (\bridge/configuration/C2340 )
    );
    defparam C19907.INIT = 16'hFFEE;
    X_LUT4 C19907(
      .ADR0 (syn177509),
      .ADR1 (syn177512),
      .ADR2 (VCC),
      .ADR3 (syn177508),
      .O (\syn177519/GROM )
    );
    defparam C19906.INIT = 16'hFEFC;
    X_LUT4 C19906(
      .ADR0 (\bridge/configuration/C2356 ),
      .ADR1 (syn120377),
      .ADR2 (syn177517),
      .ADR3 (\bridge/conf_pci_am1_out [19]),
      .O (\syn177519/FROM )
    );
    X_BUF \syn177519/YUSED (
      .I (\syn177519/GROM ),
      .O (syn177517)
    );
    X_BUF \syn177519/XUSED (
      .I (\syn177519/FROM ),
      .O (syn177519)
    );
    defparam C19936.INIT = 16'h1FFF;
    X_LUT4 C19936(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR2 (syn177397),
      .ADR3 (syn177396),
      .O (\bridge/configuration/C2356/GROM )
    );
    defparam C19935.INIT = 16'h2000;
    X_LUT4 C19935(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR2 (syn177632),
      .ADR3 (syn58393),
      .O (\bridge/configuration/C2356/FROM )
    );
    X_BUF \bridge/configuration/C2356/YUSED (
      .I (\bridge/configuration/C2356/GROM ),
      .O (syn177632)
    );
    X_BUF \bridge/configuration/C2356/XUSED (
      .I (\bridge/configuration/C2356/FROM ),
      .O (\bridge/configuration/C2356 )
    );
    defparam C19930.INIT = 16'h0080;
    X_LUT4 C19930(
      .ADR0 (syn177501),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR2 (\bridge/configuration/pci_err_data [31]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C108 ),
      .O (\syn120377/GROM )
    );
    defparam C19929.INIT = 16'h00A8;
    X_LUT4 C19929(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR1 (syn17811),
      .ADR2 (syn17815),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C116 ),
      .O (\syn120377/FROM )
    );
    X_BUF \syn120377/YUSED (
      .I (\syn120377/GROM ),
      .O (syn17815)
    );
    X_BUF \syn120377/XUSED (
      .I (\syn120377/FROM ),
      .O (syn120377)
    );
    defparam C19923.INIT = 16'h0010;
    X_LUT4 C19923(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR2 (syn60060),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .O (\syn177508/GROM )
    );
    defparam C19922.INIT = 16'h88F8;
    X_LUT4 C19922(
      .ADR0 (\bridge/configuration/C2322 ),
      .ADR1 (\bridge/conf_wb_ba1_out [19]),
      .ADR2 (syn177440),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C112 ),
      .O (\syn177508/FROM )
    );
    X_BUF \syn177508/YUSED (
      .I (\syn177508/GROM ),
      .O (syn177440)
    );
    X_BUF \syn177508/XUSED (
      .I (\syn177508/FROM ),
      .O (syn177508)
    );
    defparam C19926.INIT = 16'h0400;
    X_LUT4 C19926(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .O (\bridge/configuration/C2322/GROM )
    );
    defparam C19925.INIT = 16'h8000;
    X_LUT4 C19925(
      .ADR0 (syn177450),
      .ADR1 (syn177397),
      .ADR2 (syn177451),
      .ADR3 (syn177396),
      .O (\bridge/configuration/C2322/FROM )
    );
    X_BUF \bridge/configuration/C2322/YUSED (
      .I (\bridge/configuration/C2322/GROM ),
      .O (syn177451)
    );
    X_BUF \bridge/configuration/C2322/XUSED (
      .I (\bridge/configuration/C2322/FROM ),
      .O (\bridge/configuration/C2322 )
    );
    defparam C19918.INIT = 16'hC000;
    X_LUT4 C19918(
      .ADR0 (VCC),
      .ADR1 (syn177396),
      .ADR2 (syn177458),
      .ADR3 (syn177397),
      .O (\syn177509/GROM )
    );
    defparam C19917.INIT = 16'hF888;
    X_LUT4 C19917(
      .ADR0 (\bridge/configuration/C2302 ),
      .ADR1 (\bridge/configuration/wb_err_data [31]),
      .ADR2 (\bridge/configuration/C2292 ),
      .ADR3 (\bridge/configuration/icr_soft_res ),
      .O (\syn177509/FROM )
    );
    X_BUF \syn177509/YUSED (
      .I (\syn177509/GROM ),
      .O (\bridge/configuration/C2292 )
    );
    X_BUF \syn177509/XUSED (
      .I (\syn177509/FROM ),
      .O (syn177509)
    );
    defparam C19921.INIT = 16'h8000;
    X_LUT4 C19921(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR2 (syn58393),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .O (\bridge/configuration/C2302/GROM )
    );
    defparam C19920.INIT = 16'hC000;
    X_LUT4 C19920(
      .ADR0 (VCC),
      .ADR1 (syn177397),
      .ADR2 (syn177465),
      .ADR3 (syn177396),
      .O (\bridge/configuration/C2302/FROM )
    );
    X_BUF \bridge/configuration/C2302/YUSED (
      .I (\bridge/configuration/C2302/GROM ),
      .O (syn177465)
    );
    X_BUF \bridge/configuration/C2302/XUSED (
      .I (\bridge/configuration/C2302/FROM ),
      .O (\bridge/configuration/C2302 )
    );
    defparam C19909.INIT = 16'hC0C0;
    X_LUT4 C19909(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_pci_am1_out [19]),
      .ADR2 (\bridge/conf_pci_ba1_out [19]),
      .ADR3 (VCC),
      .O (\syn177512/GROM )
    );
    defparam C19908.INIT = 16'hFFEA;
    X_LUT4 C19908(
      .ADR0 (\bridge/configuration/C2368 ),
      .ADR1 (\bridge/configuration/C2360 ),
      .ADR2 (syn17049),
      .ADR3 (\bridge/configuration/C2320 ),
      .O (\syn177512/FROM )
    );
    X_BUF \syn177512/YUSED (
      .I (\syn177512/GROM ),
      .O (syn17049)
    );
    X_BUF \syn177512/XUSED (
      .I (\syn177512/FROM ),
      .O (syn177512)
    );
    defparam C19915.INIT = 16'h0400;
    X_LUT4 C19915(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR1 (syn177450),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR3 (syn59929),
      .O (\bridge/configuration/C2368/GROM )
    );
    defparam C19914.INIT = 16'hC000;
    X_LUT4 C19914(
      .ADR0 (VCC),
      .ADR1 (syn177396),
      .ADR2 (syn177435),
      .ADR3 (syn177397),
      .O (\bridge/configuration/C2368/FROM )
    );
    X_BUF \bridge/configuration/C2368/YUSED (
      .I (\bridge/configuration/C2368/GROM ),
      .O (syn177435)
    );
    X_BUF \bridge/configuration/C2368/XUSED (
      .I (\bridge/configuration/C2368/FROM ),
      .O (\bridge/configuration/C2368 )
    );
    defparam C19913.INIT = 16'h0020;
    X_LUT4 C19913(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR2 (syn50321),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .O (\bridge/configuration/C2360/GROM )
    );
    defparam C19912.INIT = 16'h2000;
    X_LUT4 C19912(
      .ADR0 (syn177397),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR2 (syn177446),
      .ADR3 (syn177396),
      .O (\bridge/configuration/C2360/FROM )
    );
    X_BUF \bridge/configuration/C2360/YUSED (
      .I (\bridge/configuration/C2360/GROM ),
      .O (syn177446)
    );
    X_BUF \bridge/configuration/C2360/XUSED (
      .I (\bridge/configuration/C2360/FROM ),
      .O (\bridge/configuration/C2360 )
    );
    defparam C19911.INIT = 16'h0400;
    X_LUT4 C19911(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .O (\bridge/configuration/C2320/GROM )
    );
    defparam C19910.INIT = 16'h8000;
    X_LUT4 C19910(
      .ADR0 (syn177396),
      .ADR1 (syn177397),
      .ADR2 (syn178109),
      .ADR3 (syn60060),
      .O (\bridge/configuration/C2320/FROM )
    );
    X_BUF \bridge/configuration/C2320/YUSED (
      .I (\bridge/configuration/C2320/GROM ),
      .O (syn178109)
    );
    X_BUF \bridge/configuration/C2320/XUSED (
      .I (\bridge/configuration/C2320/FROM ),
      .O (\bridge/configuration/C2320 )
    );
    defparam C19901.INIT = 16'h0020;
    X_LUT4 C19901(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR2 (syn177416),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [8]),
      .O (\syn17836/GROM )
    );
    defparam C19900.INIT = 16'h8080;
    X_LUT4 C19900(
      .ADR0 (\bridge/conf_pci_ba1_out [19]),
      .ADR1 (\bridge/conf_pci_am1_out [19]),
      .ADR2 (syn16928),
      .ADR3 (VCC),
      .O (\syn17836/FROM )
    );
    X_BUF \syn17836/YUSED (
      .I (\syn17836/GROM ),
      .O (syn16928)
    );
    X_BUF \syn17836/XUSED (
      .I (\syn17836/FROM ),
      .O (syn17836)
    );
    defparam C19952.INIT = 16'h0300;
    X_LUT4 C19952(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .O (\syn177416/GROM )
    );
    defparam C19902.INIT = 16'h2000;
    X_LUT4 C19902(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR2 (syn84030),
      .ADR3 (syn24326),
      .O (\syn177416/FROM )
    );
    X_BUF \syn177416/YUSED (
      .I (\syn177416/GROM ),
      .O (syn84030)
    );
    X_BUF \syn177416/XUSED (
      .I (\syn177416/FROM ),
      .O (syn177416)
    );
    defparam C19989.INIT = 16'h00F0;
    X_LUT4 C19989(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (N_LED),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\syn24326/GROM )
    );
    defparam C19905.INIT = 16'h0800;
    X_LUT4 C19905(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [1]),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [0]),
      .ADR2 (syn177324),
      .ADR3 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .O (\syn24326/FROM )
    );
    X_BUF \syn24326/YUSED (
      .I (\syn24326/GROM ),
      .O (syn177324)
    );
    X_BUF \syn24326/XUSED (
      .I (\syn24326/FROM ),
      .O (syn24326)
    );
    defparam C19899.INIT = 16'h2AAA;
    X_LUT4 C19899(
      .ADR0 (syn24326),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [8]),
      .ADR2 (syn177397),
      .ADR3 (syn177396),
      .O (\syn24559/GROM )
    );
    defparam C19898.INIT = 16'hA0A0;
    X_LUT4 C19898(
      .ADR0 (\bridge/configuration/C2370 ),
      .ADR1 (VCC),
      .ADR2 (syn177631),
      .ADR3 (VCC),
      .O (\syn24559/FROM )
    );
    X_BUF \syn24559/YUSED (
      .I (\syn24559/GROM ),
      .O (syn177631)
    );
    X_BUF \syn24559/XUSED (
      .I (\syn24559/FROM ),
      .O (syn24559)
    );
    defparam C19895.INIT = 16'h8000;
    X_LUT4 C19895(
      .ADR0 (syn60030),
      .ADR1 (\bridge/configuration/C3488 ),
      .ADR2 (syn59978),
      .ADR3 (syn177631),
      .O (\syn177532/GROM )
    );
    defparam C19892.INIT = 16'hEAC0;
    X_LUT4 C19892(
      .ADR0 (syn17745),
      .ADR1 (\bridge/conf_pci_ba0_out [19]),
      .ADR2 (syn16930),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [31]),
      .O (\syn177532/FROM )
    );
    X_BUF \syn177532/YUSED (
      .I (\syn177532/GROM ),
      .O (syn16930)
    );
    X_BUF \syn177532/XUSED (
      .I (\syn177532/FROM ),
      .O (syn177532)
    );
    defparam C19869.INIT = 16'hFFF8;
    X_LUT4 C19869(
      .ADR0 (syn16928),
      .ADR1 (syn17051),
      .ADR2 (syn17875),
      .ADR3 (syn16917),
      .O (\SDAT_O[30]/GROM )
    );
    defparam C19868.INIT = 16'hEEE0;
    X_LUT4 C19868(
      .ADR0 (syn177581),
      .ADR1 (syn177580),
      .ADR2 (syn177586),
      .ADR3 (syn177585),
      .O (\SDAT_O[30]/FROM )
    );
    X_BUF \SDAT_O<30>/YUSED (
      .I (\SDAT_O[30]/GROM ),
      .O (syn177586)
    );
    X_BUF \SDAT_O<30>/XUSED (
      .I (\SDAT_O[30]/FROM ),
      .O (SDAT_O[30])
    );
    defparam C19880.INIT = 16'hFF88;
    X_LUT4 C19880(
      .ADR0 (\bridge/configuration/C2304 ),
      .ADR1 (\bridge/configuration/wb_err_addr [30]),
      .ADR2 (VCC),
      .ADR3 (syn177568),
      .O (\syn177580/GROM )
    );
    defparam C19879.INIT = 16'hFFFE;
    X_LUT4 C19879(
      .ADR0 (syn177570),
      .ADR1 (syn48759),
      .ADR2 (syn177571),
      .ADR3 (syn17875),
      .O (\syn177580/FROM )
    );
    X_BUF \syn177580/YUSED (
      .I (\syn177580/GROM ),
      .O (syn177571)
    );
    X_BUF \syn177580/XUSED (
      .I (\syn177580/FROM ),
      .O (syn177580)
    );
    defparam C19883.INIT = 16'h8080;
    X_LUT4 C19883(
      .ADR0 (syn58393),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR3 (VCC),
      .O (\bridge/configuration/C2304/GROM )
    );
    defparam C19882.INIT = 16'h2000;
    X_LUT4 C19882(
      .ADR0 (syn177397),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR2 (syn177542),
      .ADR3 (syn177396),
      .O (\bridge/configuration/C2304/FROM )
    );
    X_BUF \bridge/configuration/C2304/YUSED (
      .I (\bridge/configuration/C2304/GROM ),
      .O (syn177542)
    );
    X_BUF \bridge/configuration/C2304/XUSED (
      .I (\bridge/configuration/C2304/FROM ),
      .O (\bridge/configuration/C2304 )
    );
    defparam C19876.INIT = 16'hEEEE;
    X_LUT4 C19876(
      .ADR0 (syn177569),
      .ADR1 (syn17856),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn177581/GROM )
    );
    defparam C19870.INIT = 16'hFFFE;
    X_LUT4 C19870(
      .ADR0 (syn177574),
      .ADR1 (syn177573),
      .ADR2 (syn177572),
      .ADR3 (syn177585),
      .O (\syn177581/FROM )
    );
    X_BUF \syn177581/YUSED (
      .I (\syn177581/GROM ),
      .O (syn177572)
    );
    X_BUF \syn177581/XUSED (
      .I (\syn177581/FROM ),
      .O (syn177581)
    );
    defparam C19874.INIT = 16'h0040;
    X_LUT4 C19874(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR1 (syn24500),
      .ADR2 (syn177548),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .O (\syn177573/GROM )
    );
    defparam C19873.INIT = 16'hF888;
    X_LUT4 C19873(
      .ADR0 (\bridge/configuration/C2340 ),
      .ADR1 (\bridge/configuration/pci_err_cs_bit31_24 [30]),
      .ADR2 (\bridge/configuration/C2334 ),
      .ADR3 (\bridge/configuration/pci_err_data [30]),
      .O (\syn177573/FROM )
    );
    X_BUF \syn177573/YUSED (
      .I (\syn177573/GROM ),
      .O (\bridge/configuration/C2334 )
    );
    X_BUF \syn177573/XUSED (
      .I (\syn177573/FROM ),
      .O (syn177573)
    );
    defparam C19944.INIT = 16'h8000;
    X_LUT4 C19944(
      .ADR0 (syn60043),
      .ADR1 (syn177393),
      .ADR2 (syn60044),
      .ADR3 (syn177397),
      .O (\syn16917/GROM )
    );
    defparam C19904.INIT = 16'h8080;
    X_LUT4 C19904(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [8]),
      .ADR1 (syn24326),
      .ADR2 (syn24500),
      .ADR3 (VCC),
      .O (\syn16917/FROM )
    );
    X_BUF \syn16917/YUSED (
      .I (\syn16917/GROM ),
      .O (syn24500)
    );
    X_BUF \syn16917/XUSED (
      .I (\syn16917/FROM ),
      .O (syn16917)
    );
    defparam C19854.INIT = 16'hFEFA;
    X_LUT4 C19854(
      .ADR0 (syn17912),
      .ADR1 (syn17052),
      .ADR2 (syn16917),
      .ADR3 (syn16928),
      .O (\SDAT_O[29]/GROM )
    );
    defparam C19853.INIT = 16'hFFE0;
    X_LUT4 C19853(
      .ADR0 (syn177620),
      .ADR1 (syn177616),
      .ADR2 (syn177625),
      .ADR3 (syn177624),
      .O (\SDAT_O[29]/FROM )
    );
    X_BUF \SDAT_O<29>/YUSED (
      .I (\SDAT_O[29]/GROM ),
      .O (syn177625)
    );
    X_BUF \SDAT_O<29>/XUSED (
      .I (\SDAT_O[29]/FROM ),
      .O (SDAT_O[29])
    );
    defparam C19865.INIT = 16'hFFF8;
    X_LUT4 C19865(
      .ADR0 (\bridge/configuration/wb_err_data [29]),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (syn177608),
      .ADR3 (\bridge/configuration/C2368 ),
      .O (\syn177616/GROM )
    );
    defparam C19864.INIT = 16'hFEFA;
    X_LUT4 C19864(
      .ADR0 (syn17895),
      .ADR1 (\bridge/configuration/C2304 ),
      .ADR2 (syn177611),
      .ADR3 (\bridge/configuration/wb_err_addr [29]),
      .O (\syn177616/FROM )
    );
    X_BUF \syn177616/YUSED (
      .I (\syn177616/GROM ),
      .O (syn177611)
    );
    X_BUF \syn177616/XUSED (
      .I (\syn177616/FROM ),
      .O (syn177616)
    );
    defparam C19887.INIT = 16'h0040;
    X_LUT4 C19887(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR1 (syn60060),
      .ADR2 (syn50321),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .O (\bridge/configuration/C2318/GROM )
    );
    defparam C19886.INIT = 16'h8080;
    X_LUT4 C19886(
      .ADR0 (syn177396),
      .ADR1 (syn177397),
      .ADR2 (syn177565),
      .ADR3 (VCC),
      .O (\bridge/configuration/C2318/FROM )
    );
    X_BUF \bridge/configuration/C2318/YUSED (
      .I (\bridge/configuration/C2318/GROM ),
      .O (syn177565)
    );
    X_BUF \bridge/configuration/C2318/XUSED (
      .I (\bridge/configuration/C2318/FROM ),
      .O (\bridge/configuration/C2318 )
    );
    defparam C19859.INIT = 16'hFEFA;
    X_LUT4 C19859(
      .ADR0 (syn177609),
      .ADR1 (syn16930),
      .ADR2 (syn17894),
      .ADR3 (\bridge/conf_pci_ba0_out [17]),
      .O (\syn177620/GROM )
    );
    defparam C19858.INIT = 16'hFFFA;
    X_LUT4 C19858(
      .ADR0 (syn177613),
      .ADR1 (VCC),
      .ADR2 (syn177617),
      .ADR3 (syn177614),
      .O (\syn177620/FROM )
    );
    X_BUF \syn177620/YUSED (
      .I (\syn177620/GROM ),
      .O (syn177617)
    );
    X_BUF \syn177620/XUSED (
      .I (\syn177620/FROM ),
      .O (syn177620)
    );
    defparam C19838.INIT = 16'hFFEA;
    X_LUT4 C19838(
      .ADR0 (syn177670),
      .ADR1 (\bridge/conf_pci_ba0_out [16]),
      .ADR2 (syn16930),
      .ADR3 (syn177669),
      .O (\SDAT_O[28]/GROM )
    );
    defparam C19837.INIT = 16'hFAF8;
    X_LUT4 C19837(
      .ADR0 (syn16917),
      .ADR1 (syn177665),
      .ADR2 (syn177672),
      .ADR3 (syn177664),
      .O (\SDAT_O[28]/FROM )
    );
    X_BUF \SDAT_O<28>/YUSED (
      .I (\SDAT_O[28]/GROM ),
      .O (syn177672)
    );
    X_BUF \SDAT_O<28>/XUSED (
      .I (\SDAT_O[28]/FROM ),
      .O (SDAT_O[28])
    );
    defparam C19850.INIT = 16'hECA0;
    X_LUT4 C19850(
      .ADR0 (\bridge/configuration/C2340 ),
      .ADR1 (\bridge/configuration/pci_err_data [28]),
      .ADR2 (\bridge/configuration/pci_err_cs_bit31_24 [28]),
      .ADR3 (\bridge/configuration/C2334 ),
      .O (\syn177664/GROM )
    );
    defparam C19849.INIT = 16'hFFFA;
    X_LUT4 C19849(
      .ADR0 (syn177656),
      .ADR1 (VCC),
      .ADR2 (syn177661),
      .ADR3 (syn177657),
      .O (\syn177664/FROM )
    );
    X_BUF \syn177664/YUSED (
      .I (\syn177664/GROM ),
      .O (syn177661)
    );
    X_BUF \syn177664/XUSED (
      .I (\syn177664/FROM ),
      .O (syn177664)
    );
    defparam C19844.INIT = 16'hECA0;
    X_LUT4 C19844(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [28]),
      .ADR1 (\bridge/configuration/C2356 ),
      .ADR2 (\bridge/configuration/C2354 ),
      .ADR3 (\bridge/conf_pci_am1_out [16]),
      .O (\syn177665/GROM )
    );
    defparam C19843.INIT = 16'hFFFE;
    X_LUT4 C19843(
      .ADR0 (syn177658),
      .ADR1 (syn177654),
      .ADR2 (syn177662),
      .ADR3 (syn177655),
      .O (\syn177665/FROM )
    );
    X_BUF \syn177665/YUSED (
      .I (\syn177665/GROM ),
      .O (syn177662)
    );
    X_BUF \syn177665/XUSED (
      .I (\syn177665/FROM ),
      .O (syn177665)
    );
    defparam C19841.INIT = 16'h8000;
    X_LUT4 C19841(
      .ADR0 (syn177631),
      .ADR1 (syn177632),
      .ADR2 (syn177629),
      .ADR3 (syn24500),
      .O (\syn177669/GROM )
    );
    defparam C19840.INIT = 16'hF8F0;
    X_LUT4 C19840(
      .ADR0 (\bridge/configuration/C2370 ),
      .ADR1 (syn177631),
      .ADR2 (syn17083),
      .ADR3 (\bridge/configuration/status_bit15_11 [12]),
      .O (\syn177669/FROM )
    );
    X_BUF \syn177669/YUSED (
      .I (\syn177669/GROM ),
      .O (syn17083)
    );
    X_BUF \syn177669/XUSED (
      .I (\syn177669/FROM ),
      .O (syn177669)
    );
    defparam C19822.INIT = 16'hFFFE;
    X_LUT4 C19822(
      .ADR0 (syn177701),
      .ADR1 (syn17083),
      .ADR2 (syn17990),
      .ADR3 (syn177693),
      .O (\SDAT_O[27]/GROM )
    );
    defparam C19821.INIT = 16'hFE00;
    X_LUT4 C19821(
      .ADR0 (syn177703),
      .ADR1 (syn177704),
      .ADR2 (syn177705),
      .ADR3 (syn50278),
      .O (\SDAT_O[27]/FROM )
    );
    X_BUF \SDAT_O<27>/YUSED (
      .I (\SDAT_O[27]/GROM ),
      .O (syn177705)
    );
    X_BUF \SDAT_O<27>/XUSED (
      .I (\SDAT_O[27]/FROM ),
      .O (SDAT_O[27])
    );
    defparam C19834.INIT = 16'hEAC0;
    X_LUT4 C19834(
      .ADR0 (syn17745),
      .ADR1 (\bridge/conf_pci_ba0_out [15]),
      .ADR2 (syn16930),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [27]),
      .O (\syn50278/GROM )
    );
    defparam C19833.INIT = 16'hFFFE;
    X_LUT4 C19833(
      .ADR0 (syn177710),
      .ADR1 (syn16917),
      .ADR2 (syn177711),
      .ADR3 (syn17083),
      .O (\syn50278/FROM )
    );
    X_BUF \syn50278/YUSED (
      .I (\syn50278/GROM ),
      .O (syn177711)
    );
    X_BUF \syn50278/XUSED (
      .I (\syn50278/FROM ),
      .O (syn50278)
    );
    defparam C19831.INIT = 16'hECA0;
    X_LUT4 C19831(
      .ADR0 (\bridge/configuration/C2340 ),
      .ADR1 (\bridge/configuration/C2354 ),
      .ADR2 (\bridge/configuration/pci_err_cs_bit31_24 [27]),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [27]),
      .O (\syn177703/GROM )
    );
    defparam C19830.INIT = 16'hFEFA;
    X_LUT4 C19830(
      .ADR0 (syn17971),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (syn177698),
      .ADR3 (\bridge/configuration/pci_err_data [27]),
      .O (\syn177703/FROM )
    );
    X_BUF \syn177703/YUSED (
      .I (\syn177703/GROM ),
      .O (syn177698)
    );
    X_BUF \syn177703/XUSED (
      .I (\syn177703/FROM ),
      .O (syn177703)
    );
    defparam C19829.INIT = 16'hF888;
    X_LUT4 C19829(
      .ADR0 (syn24559),
      .ADR1 (\bridge/configuration/status_bit15_11 [11]),
      .ADR2 (\bridge/configuration/C2356 ),
      .ADR3 (\bridge/conf_pci_am1_out [15]),
      .O (\syn177704/GROM )
    );
    defparam C19828.INIT = 16'hFFF8;
    X_LUT4 C19828(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [27]),
      .ADR1 (syn17745),
      .ADR2 (syn177699),
      .ADR3 (syn48759),
      .O (\syn177704/FROM )
    );
    X_BUF \syn177704/YUSED (
      .I (\syn177704/GROM ),
      .O (syn177699)
    );
    X_BUF \syn177704/XUSED (
      .I (\syn177704/FROM ),
      .O (syn177704)
    );
    defparam C19824.INIT = 16'hECA0;
    X_LUT4 C19824(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [27]),
      .ADR1 (syn17054),
      .ADR2 (\bridge/configuration/C2318 ),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn177701/GROM )
    );
    defparam C19823.INIT = 16'hFEFC;
    X_LUT4 C19823(
      .ADR0 (\bridge/configuration/C2304 ),
      .ADR1 (syn177692),
      .ADR2 (syn177694),
      .ADR3 (\bridge/configuration/wb_err_addr [27]),
      .O (\syn177701/FROM )
    );
    X_BUF \syn177701/YUSED (
      .I (\syn177701/GROM ),
      .O (syn177694)
    );
    X_BUF \syn177701/XUSED (
      .I (\syn177701/FROM ),
      .O (syn177701)
    );
    defparam C19807.INIT = 16'hFEEE;
    X_LUT4 C19807(
      .ADR0 (syn17115),
      .ADR1 (syn16917),
      .ADR2 (\bridge/conf_pci_ba0_out [14]),
      .ADR3 (syn16930),
      .O (\SDAT_O[26]/GROM )
    );
    defparam C19806.INIT = 16'hEEE0;
    X_LUT4 C19806(
      .ADR0 (syn177744),
      .ADR1 (syn177743),
      .ADR2 (syn177750),
      .ADR3 (syn177749),
      .O (\SDAT_O[26]/FROM )
    );
    X_BUF \SDAT_O<26>/YUSED (
      .I (\SDAT_O[26]/GROM ),
      .O (syn177750)
    );
    X_BUF \SDAT_O<26>/XUSED (
      .I (\SDAT_O[26]/FROM ),
      .O (SDAT_O[26])
    );
    defparam C19817.INIT = 16'hFFEC;
    X_LUT4 C19817(
      .ADR0 (\bridge/configuration/wb_err_addr [26]),
      .ADR1 (syn177732),
      .ADR2 (\bridge/configuration/C2304 ),
      .ADR3 (syn177734),
      .O (\syn177743/GROM )
    );
    defparam C19816.INIT = 16'hFEFC;
    X_LUT4 C19816(
      .ADR0 (syn17745),
      .ADR1 (syn48759),
      .ADR2 (syn177740),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [26]),
      .O (\syn177743/FROM )
    );
    X_BUF \syn177743/YUSED (
      .I (\syn177743/GROM ),
      .O (syn177740)
    );
    X_BUF \syn177743/XUSED (
      .I (\syn177743/FROM ),
      .O (syn177743)
    );
    defparam C19819.INIT = 16'hCC00;
    X_LUT4 C19819(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_pci_ba1_out [14]),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_pci_am1_out [14]),
      .O (\syn177734/GROM )
    );
    defparam C19818.INIT = 16'hEAC0;
    X_LUT4 C19818(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [26]),
      .ADR1 (\bridge/configuration/C2360 ),
      .ADR2 (syn17055),
      .ADR3 (\bridge/configuration/C2318 ),
      .O (\syn177734/FROM )
    );
    X_BUF \syn177734/YUSED (
      .I (\syn177734/GROM ),
      .O (syn17055)
    );
    X_BUF \syn177734/XUSED (
      .I (\syn177734/FROM ),
      .O (syn177734)
    );
    defparam C19811.INIT = 16'hFFEA;
    X_LUT4 C19811(
      .ADR0 (syn177733),
      .ADR1 (\bridge/conf_pci_ba0_out [14]),
      .ADR2 (syn16930),
      .ADR3 (syn18010),
      .O (\syn177744/GROM )
    );
    defparam C19810.INIT = 16'hFEFE;
    X_LUT4 C19810(
      .ADR0 (syn177738),
      .ADR1 (syn177737),
      .ADR2 (syn177741),
      .ADR3 (VCC),
      .O (\syn177744/FROM )
    );
    X_BUF \syn177744/YUSED (
      .I (\syn177744/GROM ),
      .O (syn177741)
    );
    X_BUF \syn177744/XUSED (
      .I (\syn177744/FROM ),
      .O (syn177744)
    );
    defparam C19790.INIT = 16'hFFFA;
    X_LUT4 C19790(
      .ADR0 (syn177782),
      .ADR1 (VCC),
      .ADR2 (syn177779),
      .ADR3 (syn177778),
      .O (\SDAT_O[25]/GROM )
    );
    defparam C19789.INIT = 16'hFE00;
    X_LUT4 C19789(
      .ADR0 (syn177780),
      .ADR1 (syn177781),
      .ADR2 (syn177785),
      .ADR3 (syn50276),
      .O (\SDAT_O[25]/FROM )
    );
    X_BUF \SDAT_O<25>/YUSED (
      .I (\SDAT_O[25]/GROM ),
      .O (syn177785)
    );
    X_BUF \SDAT_O<25>/XUSED (
      .I (\SDAT_O[25]/FROM ),
      .O (SDAT_O[25])
    );
    defparam C19803.INIT = 16'hFFEC;
    X_LUT4 C19803(
      .ADR0 (syn16930),
      .ADR1 (syn24559),
      .ADR2 (\bridge/conf_pci_ba0_out [13]),
      .ADR3 (syn16917),
      .O (\syn50276/GROM )
    );
    defparam C19802.INIT = 16'hFFFE;
    X_LUT4 C19802(
      .ADR0 (syn17115),
      .ADR1 (syn177790),
      .ADR2 (syn177791),
      .ADR3 (syn17083),
      .O (\syn50276/FROM )
    );
    X_BUF \syn50276/YUSED (
      .I (\syn50276/GROM ),
      .O (syn177791)
    );
    X_BUF \syn50276/XUSED (
      .I (\syn50276/FROM ),
      .O (syn50276)
    );
    defparam C19792.INIT = 16'hCC80;
    X_LUT4 C19792(
      .ADR0 (\bridge/conf_wb_ba1_out [13]),
      .ADR1 (\bridge/conf_wb_am1_out [13]),
      .ADR2 (\bridge/configuration/C2322 ),
      .ADR3 (\bridge/configuration/C2320 ),
      .O (\syn177782/GROM )
    );
    defparam C19791.INIT = 16'hFEFC;
    X_LUT4 C19791(
      .ADR0 (\bridge/conf_pci_ba0_out [13]),
      .ADR1 (syn17083),
      .ADR2 (syn18048),
      .ADR3 (syn16930),
      .O (\syn177782/FROM )
    );
    X_BUF \syn177782/YUSED (
      .I (\syn177782/GROM ),
      .O (syn18048)
    );
    X_BUF \syn177782/XUSED (
      .I (\syn177782/FROM ),
      .O (syn177782)
    );
    defparam C19775.INIT = 16'hFFEC;
    X_LUT4 C19775(
      .ADR0 (syn16928),
      .ADR1 (syn18104),
      .ADR2 (syn17057),
      .ADR3 (syn16917),
      .O (\SDAT_O[24]/GROM )
    );
    defparam C19774.INIT = 16'hFFE0;
    X_LUT4 C19774(
      .ADR0 (syn177822),
      .ADR1 (syn177826),
      .ADR2 (syn177831),
      .ADR3 (syn177830),
      .O (\SDAT_O[24]/FROM )
    );
    X_BUF \SDAT_O<24>/YUSED (
      .I (\SDAT_O[24]/GROM ),
      .O (syn177831)
    );
    X_BUF \SDAT_O<24>/XUSED (
      .I (\SDAT_O[24]/FROM ),
      .O (SDAT_O[24])
    );
    defparam C19786.INIT = 16'hFEEE;
    X_LUT4 C19786(
      .ADR0 (\bridge/configuration/C2368 ),
      .ADR1 (syn177814),
      .ADR2 (\bridge/configuration/wb_err_data [24]),
      .ADR3 (\bridge/configuration/C2302 ),
      .O (\syn177822/GROM )
    );
    defparam C19785.INIT = 16'hFEFA;
    X_LUT4 C19785(
      .ADR0 (syn18087),
      .ADR1 (\bridge/configuration/wb_err_addr [24]),
      .ADR2 (syn177817),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn177822/FROM )
    );
    X_BUF \syn177822/YUSED (
      .I (\syn177822/GROM ),
      .O (syn177817)
    );
    X_BUF \syn177822/XUSED (
      .I (\syn177822/FROM ),
      .O (syn177822)
    );
    defparam C19780.INIT = 16'hFFEC;
    X_LUT4 C19780(
      .ADR0 (syn16930),
      .ADR1 (syn177815),
      .ADR2 (\bridge/conf_pci_ba0_out [12]),
      .ADR3 (syn18086),
      .O (\syn177826/GROM )
    );
    defparam C19779.INIT = 16'hFFFC;
    X_LUT4 C19779(
      .ADR0 (VCC),
      .ADR1 (syn177819),
      .ADR2 (syn177823),
      .ADR3 (syn177820),
      .O (\syn177826/FROM )
    );
    X_BUF \syn177826/YUSED (
      .I (\syn177826/GROM ),
      .O (syn177823)
    );
    X_BUF \syn177826/XUSED (
      .I (\syn177826/FROM ),
      .O (syn177826)
    );
    defparam C19760.INIT = 16'hFFF8;
    X_LUT4 C19760(
      .ADR0 (syn17058),
      .ADR1 (syn16928),
      .ADR2 (syn17115),
      .ADR3 (syn177869),
      .O (\SDAT_O[23]/GROM )
    );
    defparam C19759.INIT = 16'hFEF0;
    X_LUT4 C19759(
      .ADR0 (syn177864),
      .ADR1 (syn177865),
      .ADR2 (syn177870),
      .ADR3 (syn16917),
      .O (\SDAT_O[23]/FROM )
    );
    X_BUF \SDAT_O<23>/YUSED (
      .I (\SDAT_O[23]/GROM ),
      .O (syn177870)
    );
    X_BUF \SDAT_O<23>/XUSED (
      .I (\SDAT_O[23]/FROM ),
      .O (SDAT_O[23])
    );
    defparam C19771.INIT = 16'hECA0;
    X_LUT4 C19771(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [23]),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (\bridge/configuration/C2354 ),
      .ADR3 (\bridge/configuration/pci_err_data [23]),
      .O (\syn177864/GROM )
    );
    defparam C19770.INIT = 16'hFFFC;
    X_LUT4 C19770(
      .ADR0 (VCC),
      .ADR1 (syn177857),
      .ADR2 (syn177861),
      .ADR3 (syn177856),
      .O (\syn177864/FROM )
    );
    X_BUF \syn177864/YUSED (
      .I (\syn177864/GROM ),
      .O (syn177861)
    );
    X_BUF \syn177864/XUSED (
      .I (\syn177864/FROM ),
      .O (syn177864)
    );
    defparam C19763.INIT = 16'hFFEA;
    X_LUT4 C19763(
      .ADR0 (syn177855),
      .ADR1 (\bridge/configuration/C2304 ),
      .ADR2 (\bridge/configuration/wb_err_addr [23]),
      .ADR3 (syn177858),
      .O (\syn177865/GROM )
    );
    defparam C19762.INIT = 16'hFEFC;
    X_LUT4 C19762(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [23]),
      .ADR1 (syn48759),
      .ADR2 (syn177863),
      .ADR3 (\bridge/configuration/C2356 ),
      .O (\syn177865/FROM )
    );
    X_BUF \syn177865/YUSED (
      .I (\syn177865/GROM ),
      .O (syn177863)
    );
    X_BUF \syn177865/XUSED (
      .I (\syn177865/FROM ),
      .O (syn177865)
    );
    defparam C19769.INIT = 16'h8888;
    X_LUT4 C19769(
      .ADR0 (\bridge/configuration/wb_addr_mask1 [23]),
      .ADR1 (\bridge/configuration/wb_base_addr1 [23]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn177855/GROM )
    );
    defparam C19768.INIT = 16'hEAC0;
    X_LUT4 C19768(
      .ADR0 (\bridge/configuration/wb_err_data [23]),
      .ADR1 (\bridge/configuration/C2322 ),
      .ADR2 (syn177838),
      .ADR3 (\bridge/configuration/C2302 ),
      .O (\syn177855/FROM )
    );
    X_BUF \syn177855/YUSED (
      .I (\syn177855/GROM ),
      .O (syn177838)
    );
    X_BUF \syn177855/XUSED (
      .I (\syn177855/FROM ),
      .O (syn177855)
    );
    defparam C19765.INIT = 16'h8888;
    X_LUT4 C19765(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [23]),
      .ADR1 (\bridge/configuration/pci_base_addr1 [23]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn177858/GROM )
    );
    defparam C19764.INIT = 16'hF888;
    X_LUT4 C19764(
      .ADR0 (\bridge/configuration/config_addr[23] ),
      .ADR1 (\bridge/configuration/C2296 ),
      .ADR2 (syn17058),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn177858/FROM )
    );
    X_BUF \syn177858/YUSED (
      .I (\syn177858/GROM ),
      .O (syn17058)
    );
    X_BUF \syn177858/XUSED (
      .I (\syn177858/FROM ),
      .O (syn177858)
    );
    defparam C19767.INIT = 16'h4040;
    X_LUT4 C19767(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR2 (syn177475),
      .ADR3 (VCC),
      .O (\bridge/configuration/C2296/GROM )
    );
    defparam C19766.INIT = 16'h4000;
    X_LUT4 C19766(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR1 (syn177396),
      .ADR2 (syn177842),
      .ADR3 (syn177397),
      .O (\bridge/configuration/C2296/FROM )
    );
    X_BUF \bridge/configuration/C2296/YUSED (
      .I (\bridge/configuration/C2296/GROM ),
      .O (syn177842)
    );
    X_BUF \bridge/configuration/C2296/XUSED (
      .I (\bridge/configuration/C2296/FROM ),
      .O (\bridge/configuration/C2296 )
    );
    defparam C19747.INIT = 16'hFCCC;
    X_LUT4 C19747(
      .ADR0 (VCC),
      .ADR1 (syn177902),
      .ADR2 (syn16930),
      .ADR3 (\bridge/configuration/pci_base_addr0 [22]),
      .O (\SDAT_O[22]/GROM )
    );
    defparam C19746.INIT = 16'hFAF8;
    X_LUT4 C19746(
      .ADR0 (syn16917),
      .ADR1 (syn177897),
      .ADR2 (syn177903),
      .ADR3 (syn177898),
      .O (\SDAT_O[22]/FROM )
    );
    X_BUF \SDAT_O<22>/YUSED (
      .I (\SDAT_O[22]/GROM ),
      .O (syn177903)
    );
    X_BUF \SDAT_O<22>/XUSED (
      .I (\SDAT_O[22]/FROM ),
      .O (SDAT_O[22])
    );
    defparam C19756.INIT = 16'hF888;
    X_LUT4 C19756(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [22]),
      .ADR1 (\bridge/configuration/C2354 ),
      .ADR2 (\bridge/configuration/C2334 ),
      .ADR3 (\bridge/configuration/pci_err_data [22]),
      .O (\syn177897/GROM )
    );
    defparam C19755.INIT = 16'hFFFA;
    X_LUT4 C19755(
      .ADR0 (syn177890),
      .ADR1 (VCC),
      .ADR2 (syn177894),
      .ADR3 (syn177889),
      .O (\syn177897/FROM )
    );
    X_BUF \syn177897/YUSED (
      .I (\syn177897/GROM ),
      .O (syn177894)
    );
    X_BUF \syn177897/XUSED (
      .I (\syn177897/FROM ),
      .O (syn177897)
    );
    defparam C19750.INIT = 16'hFEEE;
    X_LUT4 C19750(
      .ADR0 (syn177888),
      .ADR1 (syn177891),
      .ADR2 (\bridge/configuration/C2304 ),
      .ADR3 (\bridge/configuration/wb_err_addr [22]),
      .O (\syn177898/GROM )
    );
    defparam C19749.INIT = 16'hFEFC;
    X_LUT4 C19749(
      .ADR0 (\bridge/configuration/C2356 ),
      .ADR1 (syn48759),
      .ADR2 (syn177896),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [22]),
      .O (\syn177898/FROM )
    );
    X_BUF \syn177898/YUSED (
      .I (\syn177898/GROM ),
      .O (syn177896)
    );
    X_BUF \syn177898/XUSED (
      .I (\syn177898/FROM ),
      .O (syn177898)
    );
    defparam C19754.INIT = 16'hAA00;
    X_LUT4 C19754(
      .ADR0 (\bridge/configuration/wb_base_addr1 [22]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [22]),
      .O (\syn177888/GROM )
    );
    defparam C19753.INIT = 16'hF888;
    X_LUT4 C19753(
      .ADR0 (\bridge/configuration/wb_err_data [22]),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (syn177875),
      .ADR3 (\bridge/configuration/C2322 ),
      .O (\syn177888/FROM )
    );
    X_BUF \syn177888/YUSED (
      .I (\syn177888/GROM ),
      .O (syn177875)
    );
    X_BUF \syn177888/XUSED (
      .I (\syn177888/FROM ),
      .O (syn177888)
    );
    defparam C19752.INIT = 16'hAA00;
    X_LUT4 C19752(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [22]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/pci_base_addr1 [22]),
      .O (\syn177891/GROM )
    );
    defparam C19751.INIT = 16'hECA0;
    X_LUT4 C19751(
      .ADR0 (\bridge/configuration/C2360 ),
      .ADR1 (\bridge/configuration/C2296 ),
      .ADR2 (syn17059),
      .ADR3 (\bridge/configuration/config_addr[22] ),
      .O (\syn177891/FROM )
    );
    X_BUF \syn177891/YUSED (
      .I (\syn177891/GROM ),
      .O (syn17059)
    );
    X_BUF \syn177891/XUSED (
      .I (\syn177891/FROM ),
      .O (syn177891)
    );
    defparam C19741.INIT = 16'hFFFA;
    X_LUT4 C19741(
      .ADR0 (syn177927),
      .ADR1 (VCC),
      .ADR2 (syn177921),
      .ADR3 (syn177922),
      .O (\SDAT_O[21]/GROM )
    );
    defparam C19733.INIT = 16'hEEEC;
    X_LUT4 C19733(
      .ADR0 (syn16917),
      .ADR1 (syn177936),
      .ADR2 (syn177930),
      .ADR3 (syn177931),
      .O (\SDAT_O[21]/FROM )
    );
    X_BUF \SDAT_O<21>/YUSED (
      .I (\SDAT_O[21]/GROM ),
      .O (syn177930)
    );
    X_BUF \SDAT_O<21>/XUSED (
      .I (\SDAT_O[21]/FROM ),
      .O (SDAT_O[21])
    );
    defparam C19743.INIT = 16'hEAC0;
    X_LUT4 C19743(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/C2370 ),
      .ADR2 (\bridge/configuration/pci_base_addr0 [21]),
      .ADR3 (\bridge/configuration/pci_err_addr [21]),
      .O (\syn177927/GROM )
    );
    defparam C19742.INIT = 16'hFAF0;
    X_LUT4 C19742(
      .ADR0 (\bridge/configuration/C2334 ),
      .ADR1 (VCC),
      .ADR2 (syn177923),
      .ADR3 (\bridge/configuration/pci_err_data [21]),
      .O (\syn177927/FROM )
    );
    X_BUF \syn177927/YUSED (
      .I (\syn177927/GROM ),
      .O (syn177923)
    );
    X_BUF \syn177927/XUSED (
      .I (\syn177927/FROM ),
      .O (syn177927)
    );
    defparam C19737.INIT = 16'hECA0;
    X_LUT4 C19737(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [21]),
      .ADR1 (\bridge/configuration/C2354 ),
      .ADR2 (\bridge/configuration/C2356 ),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [21]),
      .O (\syn177931/GROM )
    );
    defparam C19736.INIT = 16'hFFFA;
    X_LUT4 C19736(
      .ADR0 (syn177924),
      .ADR1 (VCC),
      .ADR2 (syn177928),
      .ADR3 (syn177925),
      .O (\syn177931/FROM )
    );
    X_BUF \syn177931/YUSED (
      .I (\syn177931/GROM ),
      .O (syn177928)
    );
    X_BUF \syn177931/XUSED (
      .I (\syn177931/FROM ),
      .O (syn177931)
    );
    defparam C19735.INIT = 16'hECA0;
    X_LUT4 C19735(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [21]),
      .ADR1 (syn16928),
      .ADR2 (syn17745),
      .ADR3 (syn17060),
      .O (\syn177936/GROM )
    );
    defparam C19734.INIT = 16'hFAF0;
    X_LUT4 C19734(
      .ADR0 (\bridge/configuration/pci_base_addr0 [21]),
      .ADR1 (VCC),
      .ADR2 (syn177935),
      .ADR3 (syn16930),
      .O (\syn177936/FROM )
    );
    X_BUF \syn177936/YUSED (
      .I (\syn177936/GROM ),
      .O (syn177935)
    );
    X_BUF \syn177936/XUSED (
      .I (\syn177936/FROM ),
      .O (syn177936)
    );
    defparam C19728.INIT = 16'hFEFE;
    X_LUT4 C19728(
      .ADR0 (syn177954),
      .ADR1 (syn177955),
      .ADR2 (syn177960),
      .ADR3 (VCC),
      .O (\SDAT_O[20]/GROM )
    );
    defparam C19720.INIT = 16'hFFC8;
    X_LUT4 C19720(
      .ADR0 (syn177964),
      .ADR1 (syn16917),
      .ADR2 (syn177963),
      .ADR3 (syn177969),
      .O (\SDAT_O[20]/FROM )
    );
    X_BUF \SDAT_O<20>/YUSED (
      .I (\SDAT_O[20]/GROM ),
      .O (syn177963)
    );
    X_BUF \SDAT_O<20>/XUSED (
      .I (\SDAT_O[20]/FROM ),
      .O (SDAT_O[20])
    );
    defparam C19730.INIT = 16'hEAC0;
    X_LUT4 C19730(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/C2370 ),
      .ADR2 (\bridge/configuration/pci_base_addr0 [20]),
      .ADR3 (\bridge/configuration/pci_err_addr [20]),
      .O (\syn177960/GROM )
    );
    defparam C19729.INIT = 16'hF8F8;
    X_LUT4 C19729(
      .ADR0 (\bridge/configuration/pci_err_data [20]),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (syn177956),
      .ADR3 (VCC),
      .O (\syn177960/FROM )
    );
    X_BUF \syn177960/YUSED (
      .I (\syn177960/GROM ),
      .O (syn177956)
    );
    X_BUF \syn177960/XUSED (
      .I (\syn177960/FROM ),
      .O (syn177960)
    );
    defparam C19724.INIT = 16'hF888;
    X_LUT4 C19724(
      .ADR0 (\bridge/configuration/C2356 ),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [20]),
      .ADR2 (\bridge/configuration/C2354 ),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [20]),
      .O (\syn177964/GROM )
    );
    defparam C19723.INIT = 16'hFFFC;
    X_LUT4 C19723(
      .ADR0 (VCC),
      .ADR1 (syn177958),
      .ADR2 (syn177961),
      .ADR3 (syn177957),
      .O (\syn177964/FROM )
    );
    X_BUF \syn177964/YUSED (
      .I (\syn177964/GROM ),
      .O (syn177961)
    );
    X_BUF \syn177964/XUSED (
      .I (\syn177964/FROM ),
      .O (syn177964)
    );
    defparam C19722.INIT = 16'hF888;
    X_LUT4 C19722(
      .ADR0 (syn17745),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [20]),
      .ADR2 (syn17061),
      .ADR3 (syn16928),
      .O (\syn177969/GROM )
    );
    defparam C19721.INIT = 16'hFCF0;
    X_LUT4 C19721(
      .ADR0 (VCC),
      .ADR1 (syn16930),
      .ADR2 (syn177968),
      .ADR3 (\bridge/configuration/pci_base_addr0 [20]),
      .O (\syn177969/FROM )
    );
    X_BUF \syn177969/YUSED (
      .I (\syn177969/GROM ),
      .O (syn177968)
    );
    X_BUF \syn177969/XUSED (
      .I (\syn177969/FROM ),
      .O (syn177969)
    );
    defparam C19708.INIT = 16'hFFF8;
    X_LUT4 C19708(
      .ADR0 (syn17062),
      .ADR1 (syn16928),
      .ADR2 (syn178002),
      .ADR3 (syn17083),
      .O (\SDAT_O[19]/GROM )
    );
    defparam C19707.INIT = 16'hFEF0;
    X_LUT4 C19707(
      .ADR0 (syn177997),
      .ADR1 (syn177998),
      .ADR2 (syn178003),
      .ADR3 (syn16917),
      .O (\SDAT_O[19]/FROM )
    );
    X_BUF \SDAT_O<19>/YUSED (
      .I (\SDAT_O[19]/GROM ),
      .O (syn178003)
    );
    X_BUF \SDAT_O<19>/XUSED (
      .I (\SDAT_O[19]/FROM ),
      .O (SDAT_O[19])
    );
    defparam C19717.INIT = 16'hEAC0;
    X_LUT4 C19717(
      .ADR0 (\bridge/configuration/C2354 ),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (\bridge/configuration/pci_err_data [19]),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [19]),
      .O (\syn177997/GROM )
    );
    defparam C19716.INIT = 16'hFFFA;
    X_LUT4 C19716(
      .ADR0 (syn177989),
      .ADR1 (VCC),
      .ADR2 (syn177994),
      .ADR3 (syn177990),
      .O (\syn177997/FROM )
    );
    X_BUF \syn177997/YUSED (
      .I (\syn177997/GROM ),
      .O (syn177994)
    );
    X_BUF \syn177997/XUSED (
      .I (\syn177997/FROM ),
      .O (syn177997)
    );
    defparam C19711.INIT = 16'hFFEA;
    X_LUT4 C19711(
      .ADR0 (syn177991),
      .ADR1 (\bridge/configuration/C2304 ),
      .ADR2 (\bridge/configuration/wb_err_addr [19]),
      .ADR3 (syn177988),
      .O (\syn177998/GROM )
    );
    defparam C19710.INIT = 16'hFEFC;
    X_LUT4 C19710(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [19]),
      .ADR1 (syn48759),
      .ADR2 (syn177996),
      .ADR3 (\bridge/configuration/C2356 ),
      .O (\syn177998/FROM )
    );
    X_BUF \syn177998/YUSED (
      .I (\syn177998/GROM ),
      .O (syn177996)
    );
    X_BUF \syn177998/XUSED (
      .I (\syn177998/FROM ),
      .O (syn177998)
    );
    defparam C19715.INIT = 16'hF000;
    X_LUT4 C19715(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/wb_addr_mask1 [19]),
      .ADR3 (\bridge/configuration/wb_base_addr1 [19]),
      .O (\syn177988/GROM )
    );
    defparam C19714.INIT = 16'hEAC0;
    X_LUT4 C19714(
      .ADR0 (\bridge/configuration/C2302 ),
      .ADR1 (\bridge/configuration/C2322 ),
      .ADR2 (syn177975),
      .ADR3 (\bridge/configuration/wb_err_data [19]),
      .O (\syn177988/FROM )
    );
    X_BUF \syn177988/YUSED (
      .I (\syn177988/GROM ),
      .O (syn177975)
    );
    X_BUF \syn177988/XUSED (
      .I (\syn177988/FROM ),
      .O (syn177988)
    );
    defparam C19713.INIT = 16'hC0C0;
    X_LUT4 C19713(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [19]),
      .ADR2 (\bridge/configuration/pci_base_addr1 [19]),
      .ADR3 (VCC),
      .O (\syn177991/GROM )
    );
    defparam C19712.INIT = 16'hECA0;
    X_LUT4 C19712(
      .ADR0 (\bridge/configuration/C2360 ),
      .ADR1 (\bridge/configuration/config_addr[19] ),
      .ADR2 (syn17062),
      .ADR3 (\bridge/configuration/C2296 ),
      .O (\syn177991/FROM )
    );
    X_BUF \syn177991/YUSED (
      .I (\syn177991/GROM ),
      .O (syn17062)
    );
    X_BUF \syn177991/XUSED (
      .I (\syn177991/FROM ),
      .O (syn177991)
    );
    defparam C19695.INIT = 16'hFF88;
    X_LUT4 C19695(
      .ADR0 (\bridge/configuration/pci_base_addr0 [18]),
      .ADR1 (syn16930),
      .ADR2 (VCC),
      .ADR3 (syn178035),
      .O (\SDAT_O[18]/GROM )
    );
    defparam C19694.INIT = 16'hFCF8;
    X_LUT4 C19694(
      .ADR0 (syn178031),
      .ADR1 (syn16917),
      .ADR2 (syn178036),
      .ADR3 (syn178030),
      .O (\SDAT_O[18]/FROM )
    );
    X_BUF \SDAT_O<18>/YUSED (
      .I (\SDAT_O[18]/GROM ),
      .O (syn178036)
    );
    X_BUF \SDAT_O<18>/XUSED (
      .I (\SDAT_O[18]/FROM ),
      .O (SDAT_O[18])
    );
    defparam C19704.INIT = 16'hECA0;
    X_LUT4 C19704(
      .ADR0 (\bridge/configuration/C2354 ),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [18]),
      .ADR3 (\bridge/configuration/pci_err_data [18]),
      .O (\syn178030/GROM )
    );
    defparam C19703.INIT = 16'hFEFE;
    X_LUT4 C19703(
      .ADR0 (syn178023),
      .ADR1 (syn178022),
      .ADR2 (syn178027),
      .ADR3 (VCC),
      .O (\syn178030/FROM )
    );
    X_BUF \syn178030/YUSED (
      .I (\syn178030/GROM ),
      .O (syn178027)
    );
    X_BUF \syn178030/XUSED (
      .I (\syn178030/FROM ),
      .O (syn178030)
    );
    defparam C19698.INIT = 16'hFFEC;
    X_LUT4 C19698(
      .ADR0 (\bridge/configuration/wb_err_addr [18]),
      .ADR1 (syn178024),
      .ADR2 (\bridge/configuration/C2304 ),
      .ADR3 (syn178021),
      .O (\syn178031/GROM )
    );
    defparam C19697.INIT = 16'hFEFC;
    X_LUT4 C19697(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [18]),
      .ADR1 (syn48759),
      .ADR2 (syn178029),
      .ADR3 (\bridge/configuration/C2356 ),
      .O (\syn178031/FROM )
    );
    X_BUF \syn178031/YUSED (
      .I (\syn178031/GROM ),
      .O (syn178029)
    );
    X_BUF \syn178031/XUSED (
      .I (\syn178031/FROM ),
      .O (syn178031)
    );
    defparam C19702.INIT = 16'hCC00;
    X_LUT4 C19702(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [18]),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/wb_base_addr1 [18]),
      .O (\syn178021/GROM )
    );
    defparam C19701.INIT = 16'hECA0;
    X_LUT4 C19701(
      .ADR0 (\bridge/configuration/C2322 ),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (syn178008),
      .ADR3 (\bridge/configuration/wb_err_data [18]),
      .O (\syn178021/FROM )
    );
    X_BUF \syn178021/YUSED (
      .I (\syn178021/GROM ),
      .O (syn178008)
    );
    X_BUF \syn178021/XUSED (
      .I (\syn178021/FROM ),
      .O (syn178021)
    );
    defparam C19700.INIT = 16'hC0C0;
    X_LUT4 C19700(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_base_addr1 [18]),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [18]),
      .ADR3 (VCC),
      .O (\syn178024/GROM )
    );
    defparam C19699.INIT = 16'hECA0;
    X_LUT4 C19699(
      .ADR0 (\bridge/configuration/C2360 ),
      .ADR1 (\bridge/configuration/config_addr[18] ),
      .ADR2 (syn17063),
      .ADR3 (\bridge/configuration/C2296 ),
      .O (\syn178024/FROM )
    );
    X_BUF \syn178024/YUSED (
      .I (\syn178024/GROM ),
      .O (syn17063)
    );
    X_BUF \syn178024/XUSED (
      .I (\syn178024/FROM ),
      .O (syn178024)
    );
    defparam C19689.INIT = 16'hFEFE;
    X_LUT4 C19689(
      .ADR0 (syn178055),
      .ADR1 (syn178060),
      .ADR2 (syn178054),
      .ADR3 (VCC),
      .O (\SDAT_O[17]/GROM )
    );
    defparam C19681.INIT = 16'hFFC8;
    X_LUT4 C19681(
      .ADR0 (syn178064),
      .ADR1 (syn16917),
      .ADR2 (syn178063),
      .ADR3 (syn178069),
      .O (\SDAT_O[17]/FROM )
    );
    X_BUF \SDAT_O<17>/YUSED (
      .I (\SDAT_O[17]/GROM ),
      .O (syn178063)
    );
    X_BUF \SDAT_O<17>/XUSED (
      .I (\SDAT_O[17]/FROM ),
      .O (SDAT_O[17])
    );
    defparam C19691.INIT = 16'hEAC0;
    X_LUT4 C19691(
      .ADR0 (\bridge/configuration/pci_err_addr [17]),
      .ADR1 (\bridge/configuration/pci_base_addr0 [17]),
      .ADR2 (\bridge/configuration/C2370 ),
      .ADR3 (\bridge/configuration/C2338 ),
      .O (\syn178060/GROM )
    );
    defparam C19690.INIT = 16'hF8F8;
    X_LUT4 C19690(
      .ADR0 (\bridge/configuration/C2334 ),
      .ADR1 (\bridge/configuration/pci_err_data [17]),
      .ADR2 (syn178056),
      .ADR3 (VCC),
      .O (\syn178060/FROM )
    );
    X_BUF \syn178060/YUSED (
      .I (\syn178060/GROM ),
      .O (syn178056)
    );
    X_BUF \syn178060/XUSED (
      .I (\syn178060/FROM ),
      .O (syn178060)
    );
    defparam C19685.INIT = 16'hECA0;
    X_LUT4 C19685(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [17]),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [17]),
      .ADR2 (\bridge/configuration/C2354 ),
      .ADR3 (\bridge/configuration/C2356 ),
      .O (\syn178064/GROM )
    );
    defparam C19684.INIT = 16'hFFFA;
    X_LUT4 C19684(
      .ADR0 (syn178058),
      .ADR1 (VCC),
      .ADR2 (syn178061),
      .ADR3 (syn178057),
      .O (\syn178064/FROM )
    );
    X_BUF \syn178064/YUSED (
      .I (\syn178064/GROM ),
      .O (syn178061)
    );
    X_BUF \syn178064/XUSED (
      .I (\syn178064/FROM ),
      .O (syn178064)
    );
    defparam C19683.INIT = 16'hF888;
    X_LUT4 C19683(
      .ADR0 (syn17745),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [17]),
      .ADR2 (syn17064),
      .ADR3 (syn16928),
      .O (\syn178069/GROM )
    );
    defparam C19682.INIT = 16'hF8F8;
    X_LUT4 C19682(
      .ADR0 (\bridge/configuration/pci_base_addr0 [17]),
      .ADR1 (syn16930),
      .ADR2 (syn178068),
      .ADR3 (VCC),
      .O (\syn178069/FROM )
    );
    X_BUF \syn178069/YUSED (
      .I (\syn178069/GROM ),
      .O (syn178068)
    );
    X_BUF \syn178069/XUSED (
      .I (\syn178069/FROM ),
      .O (syn178069)
    );
    defparam C19666.INIT = 16'hFFEC;
    X_LUT4 C19666(
      .ADR0 (syn17065),
      .ADR1 (syn17118),
      .ADR2 (syn16928),
      .ADR3 (syn178106),
      .O (\SDAT_O[16]/GROM )
    );
    defparam C19665.INIT = 16'hFCF8;
    X_LUT4 C19665(
      .ADR0 (syn178102),
      .ADR1 (syn16917),
      .ADR2 (syn178107),
      .ADR3 (syn178101),
      .O (\SDAT_O[16]/FROM )
    );
    X_BUF \SDAT_O<16>/YUSED (
      .I (\SDAT_O[16]/GROM ),
      .O (syn178107)
    );
    X_BUF \SDAT_O<16>/XUSED (
      .I (\SDAT_O[16]/FROM ),
      .O (SDAT_O[16])
    );
    defparam C19677.INIT = 16'hEEAA;
    X_LUT4 C19677(
      .ADR0 (syn178094),
      .ADR1 (\bridge/configuration/pci_err_data [16]),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C2334 ),
      .O (\syn178101/GROM )
    );
    defparam C19676.INIT = 16'hFEFE;
    X_LUT4 C19676(
      .ADR0 (syn178093),
      .ADR1 (syn178092),
      .ADR2 (syn178098),
      .ADR3 (VCC),
      .O (\syn178101/FROM )
    );
    X_BUF \syn178101/YUSED (
      .I (\syn178101/GROM ),
      .O (syn178098)
    );
    X_BUF \syn178101/XUSED (
      .I (\syn178101/FROM ),
      .O (syn178101)
    );
    defparam C19672.INIT = 16'hF888;
    X_LUT4 C19672(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [16]),
      .ADR1 (\bridge/configuration/C2356 ),
      .ADR2 (\bridge/configuration/C2354 ),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [16]),
      .O (\syn178102/GROM )
    );
    defparam C19671.INIT = 16'hFFFC;
    X_LUT4 C19671(
      .ADR0 (VCC),
      .ADR1 (syn178095),
      .ADR2 (syn178099),
      .ADR3 (syn178096),
      .O (\syn178102/FROM )
    );
    X_BUF \syn178102/YUSED (
      .I (\syn178102/GROM ),
      .O (syn178099)
    );
    X_BUF \syn178102/XUSED (
      .I (\syn178102/FROM ),
      .O (syn178102)
    );
    defparam C19924.INIT = 16'h0011;
    X_LUT4 C19924(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .O (\syn17772/GROM )
    );
    defparam C19669.INIT = 16'h73FF;
    X_LUT4 C19669(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR1 (syn177396),
      .ADR2 (syn178071),
      .ADR3 (syn177397),
      .O (\syn17772/FROM )
    );
    X_BUF \syn17772/YUSED (
      .I (\syn17772/GROM ),
      .O (syn178071)
    );
    X_BUF \syn17772/XUSED (
      .I (\syn17772/FROM ),
      .O (syn17772)
    );
    defparam C19651.INIT = 16'hFFF8;
    X_LUT4 C19651(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [15]),
      .ADR1 (syn17745),
      .ADR2 (syn18431),
      .ADR3 (syn178144),
      .O (\SDAT_O[15]/GROM )
    );
    defparam C19650.INIT = 16'hFEF0;
    X_LUT4 C19650(
      .ADR0 (syn178140),
      .ADR1 (syn178139),
      .ADR2 (syn178145),
      .ADR3 (syn16917),
      .O (\SDAT_O[15]/FROM )
    );
    X_BUF \SDAT_O<15>/YUSED (
      .I (\SDAT_O[15]/GROM ),
      .O (syn178145)
    );
    X_BUF \SDAT_O<15>/XUSED (
      .I (\SDAT_O[15]/FROM ),
      .O (SDAT_O[15])
    );
    defparam C19662.INIT = 16'hECA0;
    X_LUT4 C19662(
      .ADR0 (\bridge/configuration/C2334 ),
      .ADR1 (\bridge/configuration/pci_tran_addr1 [15]),
      .ADR2 (\bridge/configuration/pci_err_data [15]),
      .ADR3 (\bridge/configuration/C2354 ),
      .O (\syn178139/GROM )
    );
    defparam C19661.INIT = 16'hFFFC;
    X_LUT4 C19661(
      .ADR0 (VCC),
      .ADR1 (syn178132),
      .ADR2 (syn178136),
      .ADR3 (syn178131),
      .O (\syn178139/FROM )
    );
    X_BUF \syn178139/YUSED (
      .I (\syn178139/GROM ),
      .O (syn178136)
    );
    X_BUF \syn178139/XUSED (
      .I (\syn178139/FROM ),
      .O (syn178139)
    );
    defparam C19656.INIT = 16'hFFEA;
    X_LUT4 C19656(
      .ADR0 (syn178133),
      .ADR1 (\bridge/configuration/C2304 ),
      .ADR2 (\bridge/configuration/wb_err_addr [15]),
      .ADR3 (syn178130),
      .O (\syn178140/GROM )
    );
    defparam C19655.INIT = 16'hFFF8;
    X_LUT4 C19655(
      .ADR0 (\bridge/configuration/C2356 ),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [15]),
      .ADR2 (syn178138),
      .ADR3 (syn48759),
      .O (\syn178140/FROM )
    );
    X_BUF \syn178140/YUSED (
      .I (\syn178140/GROM ),
      .O (syn178138)
    );
    X_BUF \syn178140/XUSED (
      .I (\syn178140/FROM ),
      .O (syn178140)
    );
    defparam C19660.INIT = 16'hAA00;
    X_LUT4 C19660(
      .ADR0 (\bridge/configuration/wb_addr_mask1 [15]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/wb_base_addr1 [15]),
      .O (\syn178130/GROM )
    );
    defparam C19659.INIT = 16'hF888;
    X_LUT4 C19659(
      .ADR0 (\bridge/configuration/wb_err_data [15]),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (syn178117),
      .ADR3 (\bridge/configuration/C2322 ),
      .O (\syn178130/FROM )
    );
    X_BUF \syn178130/YUSED (
      .I (\syn178130/GROM ),
      .O (syn178117)
    );
    X_BUF \syn178130/XUSED (
      .I (\syn178130/FROM ),
      .O (syn178130)
    );
    defparam C19658.INIT = 16'hC0C0;
    X_LUT4 C19658(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_base_addr1 [15]),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [15]),
      .ADR3 (VCC),
      .O (\syn178133/GROM )
    );
    defparam C19657.INIT = 16'hF888;
    X_LUT4 C19657(
      .ADR0 (\bridge/configuration/config_addr[15] ),
      .ADR1 (\bridge/configuration/C2296 ),
      .ADR2 (syn17066),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn178133/FROM )
    );
    X_BUF \syn178133/YUSED (
      .I (\syn178133/GROM ),
      .O (syn17066)
    );
    X_BUF \syn178133/XUSED (
      .I (\syn178133/FROM ),
      .O (syn178133)
    );
    defparam C19653.INIT = 16'h8000;
    X_LUT4 C19653(
      .ADR0 (syn178109),
      .ADR1 (syn24500),
      .ADR2 (syn177632),
      .ADR3 (syn177631),
      .O (\syn178144/GROM )
    );
    defparam C19652.INIT = 16'hECA0;
    X_LUT4 C19652(
      .ADR0 (\bridge/conf_latency_tim_out [7]),
      .ADR1 (syn16930),
      .ADR2 (syn17067),
      .ADR3 (\bridge/configuration/pci_base_addr0 [15]),
      .O (\syn178144/FROM )
    );
    X_BUF \syn178144/YUSED (
      .I (\syn178144/GROM ),
      .O (syn17067)
    );
    X_BUF \syn178144/XUSED (
      .I (\syn178144/FROM ),
      .O (syn178144)
    );
    defparam C19637.INIT = 16'hFEFC;
    X_LUT4 C19637(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [14]),
      .ADR1 (syn18468),
      .ADR2 (syn178179),
      .ADR3 (syn17745),
      .O (\SDAT_O[14]/GROM )
    );
    defparam C19636.INIT = 16'hFCF8;
    X_LUT4 C19636(
      .ADR0 (syn178174),
      .ADR1 (syn16917),
      .ADR2 (syn178180),
      .ADR3 (syn178175),
      .O (\SDAT_O[14]/FROM )
    );
    X_BUF \SDAT_O<14>/YUSED (
      .I (\SDAT_O[14]/GROM ),
      .O (syn178180)
    );
    X_BUF \SDAT_O<14>/XUSED (
      .I (\SDAT_O[14]/FROM ),
      .O (SDAT_O[14])
    );
    defparam C19647.INIT = 16'hF888;
    X_LUT4 C19647(
      .ADR0 (\bridge/configuration/C2334 ),
      .ADR1 (\bridge/configuration/pci_err_data [14]),
      .ADR2 (\bridge/configuration/C2354 ),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [14]),
      .O (\syn178174/GROM )
    );
    defparam C19646.INIT = 16'hFFFC;
    X_LUT4 C19646(
      .ADR0 (VCC),
      .ADR1 (syn178166),
      .ADR2 (syn178171),
      .ADR3 (syn178167),
      .O (\syn178174/FROM )
    );
    X_BUF \syn178174/YUSED (
      .I (\syn178174/GROM ),
      .O (syn178171)
    );
    X_BUF \syn178174/XUSED (
      .I (\syn178174/FROM ),
      .O (syn178174)
    );
    defparam C19641.INIT = 16'hFEEE;
    X_LUT4 C19641(
      .ADR0 (syn178165),
      .ADR1 (syn178168),
      .ADR2 (\bridge/configuration/C2304 ),
      .ADR3 (\bridge/configuration/wb_err_addr [14]),
      .O (\syn178175/GROM )
    );
    defparam C19640.INIT = 16'hFFF8;
    X_LUT4 C19640(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [14]),
      .ADR1 (\bridge/configuration/C2356 ),
      .ADR2 (syn178173),
      .ADR3 (syn48759),
      .O (\syn178175/FROM )
    );
    X_BUF \syn178175/YUSED (
      .I (\syn178175/GROM ),
      .O (syn178173)
    );
    X_BUF \syn178175/XUSED (
      .I (\syn178175/FROM ),
      .O (syn178175)
    );
    defparam C19645.INIT = 16'hAA00;
    X_LUT4 C19645(
      .ADR0 (\bridge/configuration/wb_base_addr1 [14]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [14]),
      .O (\syn178165/GROM )
    );
    defparam C19644.INIT = 16'hF888;
    X_LUT4 C19644(
      .ADR0 (\bridge/configuration/C2302 ),
      .ADR1 (\bridge/configuration/wb_err_data [14]),
      .ADR2 (syn178152),
      .ADR3 (\bridge/configuration/C2322 ),
      .O (\syn178165/FROM )
    );
    X_BUF \syn178165/YUSED (
      .I (\syn178165/GROM ),
      .O (syn178152)
    );
    X_BUF \syn178165/XUSED (
      .I (\syn178165/FROM ),
      .O (syn178165)
    );
    defparam C19643.INIT = 16'hAA00;
    X_LUT4 C19643(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [14]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/pci_base_addr1 [14]),
      .O (\syn178168/GROM )
    );
    defparam C19642.INIT = 16'hEAC0;
    X_LUT4 C19642(
      .ADR0 (\bridge/configuration/config_addr[14] ),
      .ADR1 (\bridge/configuration/C2360 ),
      .ADR2 (syn17068),
      .ADR3 (\bridge/configuration/C2296 ),
      .O (\syn178168/FROM )
    );
    X_BUF \syn178168/YUSED (
      .I (\syn178168/GROM ),
      .O (syn17068)
    );
    X_BUF \syn178168/XUSED (
      .I (\syn178168/FROM ),
      .O (syn178168)
    );
    defparam C19623.INIT = 16'hFFF8;
    X_LUT4 C19623(
      .ADR0 (\bridge/configuration/pci_base_addr0 [13]),
      .ADR1 (syn16930),
      .ADR2 (syn178214),
      .ADR3 (syn178213),
      .O (\SDAT_O[13]/GROM )
    );
    defparam C19622.INIT = 16'hFCF0;
    X_LUT4 C19622(
      .ADR0 (VCC),
      .ADR1 (syn18511),
      .ADR2 (syn178216),
      .ADR3 (syn16917),
      .O (\SDAT_O[13]/FROM )
    );
    X_BUF \SDAT_O<13>/YUSED (
      .I (\SDAT_O[13]/GROM ),
      .O (syn178216)
    );
    X_BUF \SDAT_O<13>/XUSED (
      .I (\SDAT_O[13]/FROM ),
      .O (SDAT_O[13])
    );
    defparam C19633.INIT = 16'hEEEE;
    X_LUT4 C19633(
      .ADR0 (syn178200),
      .ADR1 (syn178201),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn18511/GROM )
    );
    defparam C19626.INIT = 16'hFFFE;
    X_LUT4 C19626(
      .ADR0 (syn178207),
      .ADR1 (syn178208),
      .ADR2 (syn178205),
      .ADR3 (syn178206),
      .O (\syn18511/FROM )
    );
    X_BUF \syn18511/YUSED (
      .I (\syn18511/GROM ),
      .O (syn178205)
    );
    X_BUF \syn18511/XUSED (
      .I (\syn18511/FROM ),
      .O (syn18511)
    );
    defparam C19632.INIT = 16'hEAC0;
    X_LUT4 C19632(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/C2370 ),
      .ADR2 (\bridge/configuration/pci_base_addr0 [13]),
      .ADR3 (\bridge/configuration/pci_err_addr [13]),
      .O (\syn178206/GROM )
    );
    defparam C19631.INIT = 16'hF8F8;
    X_LUT4 C19631(
      .ADR0 (\bridge/configuration/pci_err_data [13]),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (syn178202),
      .ADR3 (VCC),
      .O (\syn178206/FROM )
    );
    X_BUF \syn178206/YUSED (
      .I (\syn178206/GROM ),
      .O (syn178202)
    );
    X_BUF \syn178206/XUSED (
      .I (\syn178206/FROM ),
      .O (syn178206)
    );
    defparam C19628.INIT = 16'hEAC0;
    X_LUT4 C19628(
      .ADR0 (\bridge/configuration/C2304 ),
      .ADR1 (\bridge/configuration/config_addr[13] ),
      .ADR2 (\bridge/configuration/C2296 ),
      .ADR3 (\bridge/configuration/wb_err_addr [13]),
      .O (\syn178208/GROM )
    );
    defparam C19627.INIT = 16'hFFF8;
    X_LUT4 C19627(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [13]),
      .ADR2 (syn178204),
      .ADR3 (syn18491),
      .O (\syn178208/FROM )
    );
    X_BUF \syn178208/YUSED (
      .I (\syn178208/GROM ),
      .O (syn178204)
    );
    X_BUF \syn178208/XUSED (
      .I (\syn178208/FROM ),
      .O (syn178208)
    );
    defparam C19668.INIT = 16'h2000;
    X_LUT4 C19668(
      .ADR0 (syn17772),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR2 (syn24326),
      .ADR3 (syn177632),
      .O (\syn178213/GROM )
    );
    defparam C19625.INIT = 16'hF8F0;
    X_LUT4 C19625(
      .ADR0 (\bridge/configuration/pci_base_addr1 [13]),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [13]),
      .ADR2 (syn17118),
      .ADR3 (syn16928),
      .O (\syn178213/FROM )
    );
    X_BUF \syn178213/YUSED (
      .I (\syn178213/GROM ),
      .O (syn17118)
    );
    X_BUF \syn178213/XUSED (
      .I (\syn178213/FROM ),
      .O (syn178213)
    );
    defparam C19609.INIT = 16'hFFEA;
    X_LUT4 C19609(
      .ADR0 (syn18543),
      .ADR1 (syn17745),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [12]),
      .ADR3 (syn178250),
      .O (\SDAT_O[12]/GROM )
    );
    defparam C19608.INIT = 16'hFEF0;
    X_LUT4 C19608(
      .ADR0 (syn178245),
      .ADR1 (syn178246),
      .ADR2 (syn178251),
      .ADR3 (syn16917),
      .O (\SDAT_O[12]/FROM )
    );
    X_BUF \SDAT_O<12>/YUSED (
      .I (\SDAT_O[12]/GROM ),
      .O (syn178251)
    );
    X_BUF \SDAT_O<12>/XUSED (
      .I (\SDAT_O[12]/FROM ),
      .O (SDAT_O[12])
    );
    defparam C19618.INIT = 16'hECEC;
    X_LUT4 C19618(
      .ADR0 (\bridge/configuration/pci_err_data [12]),
      .ADR1 (syn178238),
      .ADR2 (\bridge/configuration/C2334 ),
      .ADR3 (VCC),
      .O (\syn178245/GROM )
    );
    defparam C19617.INIT = 16'hFEFE;
    X_LUT4 C19617(
      .ADR0 (syn178237),
      .ADR1 (syn178236),
      .ADR2 (syn178242),
      .ADR3 (VCC),
      .O (\syn178245/FROM )
    );
    X_BUF \syn178245/YUSED (
      .I (\syn178245/GROM ),
      .O (syn178242)
    );
    X_BUF \syn178245/XUSED (
      .I (\syn178245/FROM ),
      .O (syn178245)
    );
    defparam C19613.INIT = 16'hECA0;
    X_LUT4 C19613(
      .ADR0 (\bridge/configuration/C2354 ),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [12]),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [12]),
      .ADR3 (\bridge/configuration/C2356 ),
      .O (\syn178246/GROM )
    );
    defparam C19612.INIT = 16'hFFFA;
    X_LUT4 C19612(
      .ADR0 (syn178239),
      .ADR1 (VCC),
      .ADR2 (syn178243),
      .ADR3 (syn178240),
      .O (\syn178246/FROM )
    );
    X_BUF \syn178246/YUSED (
      .I (\syn178246/GROM ),
      .O (syn178243)
    );
    X_BUF \syn178246/XUSED (
      .I (\syn178246/FROM ),
      .O (syn178246)
    );
    defparam C19599.INIT = 16'hEAC0;
    X_LUT4 C19599(
      .ADR0 (syn17067),
      .ADR1 (syn17072),
      .ADR2 (\bridge/configuration/pci_err_data [11]),
      .ADR3 (\bridge/conf_latency_tim_out [3]),
      .O (\SDAT_O[11]/GROM )
    );
    defparam C19598.INIT = 16'hFFFE;
    X_LUT4 C19598(
      .ADR0 (syn178266),
      .ADR1 (syn178265),
      .ADR2 (syn178268),
      .ADR3 (syn18567),
      .O (\SDAT_O[11]/FROM )
    );
    X_BUF \SDAT_O<11>/YUSED (
      .I (\SDAT_O[11]/GROM ),
      .O (syn178268)
    );
    X_BUF \SDAT_O<11>/XUSED (
      .I (\SDAT_O[11]/FROM ),
      .O (SDAT_O[11])
    );
    defparam C19605.INIT = 16'hF000;
    X_LUT4 C19605(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/C2302 ),
      .ADR3 (syn16917),
      .O (\syn178265/GROM )
    );
    defparam C19604.INIT = 16'hEAC0;
    X_LUT4 C19604(
      .ADR0 (\bridge/configuration/pci_err_addr [11]),
      .ADR1 (\bridge/configuration/wb_err_data [11]),
      .ADR2 (syn17075),
      .ADR3 (syn17071),
      .O (\syn178265/FROM )
    );
    X_BUF \syn178265/YUSED (
      .I (\syn178265/GROM ),
      .O (syn17075)
    );
    X_BUF \syn178265/XUSED (
      .I (\syn178265/FROM ),
      .O (syn178265)
    );
    defparam C19602.INIT = 16'hA0A0;
    X_LUT4 C19602(
      .ADR0 (syn16917),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/C2296 ),
      .ADR3 (VCC),
      .O (\syn178266/GROM )
    );
    defparam C19601.INIT = 16'hEAC0;
    X_LUT4 C19601(
      .ADR0 (syn17073),
      .ADR1 (\bridge/configuration/config_addr[11] ),
      .ADR2 (syn17076),
      .ADR3 (\bridge/configuration/wb_err_addr [11]),
      .O (\syn178266/FROM )
    );
    X_BUF \syn178266/YUSED (
      .I (\syn178266/GROM ),
      .O (syn17076)
    );
    X_BUF \syn178266/XUSED (
      .I (\syn178266/FROM ),
      .O (syn178266)
    );
    defparam C19583.INIT = 16'hFEFC;
    X_LUT4 C19583(
      .ADR0 (syn16984),
      .ADR1 (syn178292),
      .ADR2 (syn18585),
      .ADR3 (\bridge/configuration/pci_err_addr [10]),
      .O (\SDAT_O[10]/GROM )
    );
    defparam C19582.INIT = 16'hFE00;
    X_LUT4 C19582(
      .ADR0 (syn178294),
      .ADR1 (syn178293),
      .ADR2 (syn178295),
      .ADR3 (syn24466),
      .O (\SDAT_O[10]/FROM )
    );
    X_BUF \SDAT_O<10>/YUSED (
      .I (\SDAT_O[10]/GROM ),
      .O (syn178295)
    );
    X_BUF \SDAT_O<10>/XUSED (
      .I (\SDAT_O[10]/FROM ),
      .O (SDAT_O[10])
    );
    defparam C19590.INIT = 16'hA000;
    X_LUT4 C19590(
      .ADR0 (syn16936),
      .ADR1 (VCC),
      .ADR2 (syn178109),
      .ADR3 (syn24500),
      .O (\syn178294/GROM )
    );
    defparam C19589.INIT = 16'hEAC0;
    X_LUT4 C19589(
      .ADR0 (\bridge/configuration/pci_err_data [10]),
      .ADR1 (\bridge/conf_latency_tim_out [2]),
      .ADR2 (syn17081),
      .ADR3 (syn17077),
      .O (\syn178294/FROM )
    );
    X_BUF \syn178294/YUSED (
      .I (\syn178294/GROM ),
      .O (syn17081)
    );
    X_BUF \syn178294/XUSED (
      .I (\syn178294/FROM ),
      .O (syn178294)
    );
    defparam C19896.INIT = 16'h3FFF;
    X_LUT4 C19896(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR2 (syn177396),
      .ADR3 (syn177397),
      .O (\syn16936/GROM )
    );
    defparam C19591.INIT = 16'h00A0;
    X_LUT4 C19591(
      .ADR0 (syn59978),
      .ADR1 (VCC),
      .ADR2 (syn60030),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .O (\syn16936/FROM )
    );
    X_BUF \syn16936/YUSED (
      .I (\syn16936/GROM ),
      .O (syn60030)
    );
    X_BUF \syn16936/XUSED (
      .I (\syn16936/FROM ),
      .O (syn16936)
    );
    defparam C19585.INIT = 16'hC0C0;
    X_LUT4 C19585(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR2 (\bridge/configuration/C2296 ),
      .ADR3 (VCC),
      .O (\syn178292/GROM )
    );
    defparam C19584.INIT = 16'hF888;
    X_LUT4 C19584(
      .ADR0 (syn17078),
      .ADR1 (\bridge/configuration/wb_err_addr [10]),
      .ADR2 (syn17079),
      .ADR3 (\bridge/configuration/config_addr[10] ),
      .O (\syn178292/FROM )
    );
    X_BUF \syn178292/YUSED (
      .I (\syn178292/GROM ),
      .O (syn17079)
    );
    X_BUF \syn178292/XUSED (
      .I (\syn178292/FROM ),
      .O (syn178292)
    );
    defparam C19575.INIT = 16'hFEEE;
    X_LUT4 C19575(
      .ADR0 (syn17119),
      .ADR1 (syn178311),
      .ADR2 (\bridge/configuration/pci_err_addr [9]),
      .ADR3 (syn16984),
      .O (\SDAT_O[9]/GROM )
    );
    defparam C19574.INIT = 16'hCCC8;
    X_LUT4 C19574(
      .ADR0 (syn178313),
      .ADR1 (syn24468),
      .ADR2 (syn178314),
      .ADR3 (syn178312),
      .O (\SDAT_O[9]/FROM )
    );
    X_BUF \SDAT_O<9>/YUSED (
      .I (\SDAT_O[9]/GROM ),
      .O (syn178314)
    );
    X_BUF \SDAT_O<9>/XUSED (
      .I (\SDAT_O[9]/FROM ),
      .O (SDAT_O[9])
    );
    defparam C19580.INIT = 16'hECA0;
    X_LUT4 C19580(
      .ADR0 (syn17080),
      .ADR1 (syn17074),
      .ADR2 (\bridge/configuration/wb_err_cs_bit10_8 [9]),
      .ADR3 (\bridge/configuration/wb_err_data [9]),
      .O (\syn178312/GROM )
    );
    defparam C19579.INIT = 16'hF8F8;
    X_LUT4 C19579(
      .ADR0 (syn17745),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [9]),
      .ADR2 (syn178309),
      .ADR3 (VCC),
      .O (\syn178312/FROM )
    );
    X_BUF \syn178312/YUSED (
      .I (\syn178312/GROM ),
      .O (syn178309)
    );
    X_BUF \syn178312/XUSED (
      .I (\syn178312/FROM ),
      .O (syn178312)
    );
    defparam C19562.INIT = 16'hFEFA;
    X_LUT4 C19562(
      .ADR0 (syn178338),
      .ADR1 (syn17745),
      .ADR2 (syn178334),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [8]),
      .O (\SDAT_O[8]/GROM )
    );
    defparam C19561.INIT = 16'hFE00;
    X_LUT4 C19561(
      .ADR0 (syn178341),
      .ADR1 (syn178340),
      .ADR2 (syn178342),
      .ADR3 (syn24470),
      .O (\SDAT_O[8]/FROM )
    );
    X_BUF \SDAT_O<8>/YUSED (
      .I (\SDAT_O[8]/GROM ),
      .O (syn178342)
    );
    X_BUF \SDAT_O<8>/XUSED (
      .I (\SDAT_O[8]/FROM ),
      .O (SDAT_O[8])
    );
    defparam C19571.INIT = 16'hECCC;
    X_LUT4 C19571(
      .ADR0 (\bridge/configuration/wb_err_addr [8]),
      .ADR1 (syn18636),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn178340/GROM )
    );
    defparam C19570.INIT = 16'hFAF0;
    X_LUT4 C19570(
      .ADR0 (syn17081),
      .ADR1 (VCC),
      .ADR2 (syn178335),
      .ADR3 (\bridge/conf_latency_tim_out [0]),
      .O (\syn178340/FROM )
    );
    X_BUF \syn178340/YUSED (
      .I (\syn178340/GROM ),
      .O (syn178335)
    );
    X_BUF \syn178340/XUSED (
      .I (\syn178340/FROM ),
      .O (syn178340)
    );
    defparam C19568.INIT = 16'hECCC;
    X_LUT4 C19568(
      .ADR0 (\bridge/configuration/C2340 ),
      .ADR1 (syn17119),
      .ADR2 (\bridge/conf_pci_err_pending_out ),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .O (\syn178341/GROM )
    );
    defparam C19567.INIT = 16'hFEFA;
    X_LUT4 C19567(
      .ADR0 (syn17084),
      .ADR1 (\bridge/configuration/pci_err_addr [8]),
      .ADR2 (syn178337),
      .ADR3 (syn16984),
      .O (\syn178341/FROM )
    );
    X_BUF \syn178341/YUSED (
      .I (\syn178341/GROM ),
      .O (syn178337)
    );
    X_BUF \syn178341/XUSED (
      .I (\syn178341/FROM ),
      .O (syn178341)
    );
    defparam C19566.INIT = 16'h8800;
    X_LUT4 C19566(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR1 (\bridge/conf_wb_err_pending_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C2308 ),
      .O (\syn178334/GROM )
    );
    defparam C19565.INIT = 16'hF0F8;
    X_LUT4 C19565(
      .ADR0 (\bridge/conf_serr_enable_out ),
      .ADR1 (\bridge/configuration/C2370 ),
      .ADR2 (syn18632),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .O (\syn178334/FROM )
    );
    X_BUF \syn178334/YUSED (
      .I (\syn178334/GROM ),
      .O (syn18632)
    );
    X_BUF \syn178334/XUSED (
      .I (\syn178334/FROM ),
      .O (syn178334)
    );
    defparam C19564.INIT = 16'hA000;
    X_LUT4 C19564(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/C2296 ),
      .ADR3 (\bridge/configuration/config_addr[8] ),
      .O (\syn178338/GROM )
    );
    defparam C19563.INIT = 16'hF8F0;
    X_LUT4 C19563(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR1 (\bridge/configuration/pci_err_data [8]),
      .ADR2 (syn18633),
      .ADR3 (\bridge/configuration/C2334 ),
      .O (\syn178338/FROM )
    );
    X_BUF \syn178338/YUSED (
      .I (\syn178338/GROM ),
      .O (syn18633)
    );
    X_BUF \syn178338/XUSED (
      .I (\syn178338/FROM ),
      .O (syn178338)
    );
    defparam C19555.INIT = 16'hF888;
    X_LUT4 C19555(
      .ADR0 (syn17072),
      .ADR1 (\bridge/configuration/pci_err_data [7]),
      .ADR2 (syn17083),
      .ADR3 (\bridge/configuration/interrupt_line [7]),
      .O (\SDAT_O[7]/GROM )
    );
    defparam C19554.INIT = 16'hFFFE;
    X_LUT4 C19554(
      .ADR0 (syn18659),
      .ADR1 (syn178356),
      .ADR2 (syn178358),
      .ADR3 (syn178357),
      .O (\SDAT_O[7]/FROM )
    );
    X_BUF \SDAT_O<7>/YUSED (
      .I (\SDAT_O[7]/GROM ),
      .O (syn178358)
    );
    X_BUF \SDAT_O<7>/XUSED (
      .I (\SDAT_O[7]/FROM ),
      .O (SDAT_O[7])
    );
    defparam C19557.INIT = 16'h8080;
    X_LUT4 C19557(
      .ADR0 (\bridge/configuration/pci_err_addr [7]),
      .ADR1 (\bridge/configuration/C2338 ),
      .ADR2 (syn16917),
      .ADR3 (VCC),
      .O (\syn178357/GROM )
    );
    defparam C19556.INIT = 16'hFFF8;
    X_LUT4 C19556(
      .ADR0 (syn17745),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [7]),
      .ADR2 (syn18658),
      .ADR3 (syn18655),
      .O (\syn178357/FROM )
    );
    X_BUF \syn178357/YUSED (
      .I (\syn178357/GROM ),
      .O (syn18658)
    );
    X_BUF \syn178357/XUSED (
      .I (\syn178357/FROM ),
      .O (syn178357)
    );
    defparam C19546.INIT = 16'hFFEC;
    X_LUT4 C19546(
      .ADR0 (syn17078),
      .ADR1 (syn178373),
      .ADR2 (\bridge/configuration/wb_err_addr [6]),
      .ADR3 (syn18681),
      .O (\SDAT_O[6]/GROM )
    );
    defparam C19545.INIT = 16'hAAA8;
    X_LUT4 C19545(
      .ADR0 (syn24472),
      .ADR1 (syn178376),
      .ADR2 (syn178377),
      .ADR3 (syn178375),
      .O (\SDAT_O[6]/FROM )
    );
    X_BUF \SDAT_O<6>/YUSED (
      .I (\SDAT_O[6]/GROM ),
      .O (syn178377)
    );
    X_BUF \SDAT_O<6>/XUSED (
      .I (\SDAT_O[6]/FROM ),
      .O (SDAT_O[6])
    );
    defparam C19551.INIT = 16'hF8F0;
    X_LUT4 C19551(
      .ADR0 (\bridge/configuration/C2302 ),
      .ADR1 (\bridge/configuration/wb_err_data [6]),
      .ADR2 (syn18670),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .O (\syn178375/GROM )
    );
    defparam C19550.INIT = 16'hFCF0;
    X_LUT4 C19550(
      .ADR0 (VCC),
      .ADR1 (syn17084),
      .ADR2 (syn178372),
      .ADR3 (\bridge/configuration/interrupt_line [6]),
      .O (\syn178375/FROM )
    );
    X_BUF \syn178375/YUSED (
      .I (\syn178375/GROM ),
      .O (syn178372)
    );
    X_BUF \syn178375/XUSED (
      .I (\syn178375/FROM ),
      .O (syn178375)
    );
    defparam C19539.INIT = 16'hFFEC;
    X_LUT4 C19539(
      .ADR0 (\bridge/configuration/config_addr[5] ),
      .ADR1 (syn17119),
      .ADR2 (syn17079),
      .ADR3 (syn178392),
      .O (\SDAT_O[5]/GROM )
    );
    defparam C19538.INIT = 16'hFE00;
    X_LUT4 C19538(
      .ADR0 (syn178393),
      .ADR1 (syn178394),
      .ADR2 (syn178395),
      .ADR3 (syn24474),
      .O (\SDAT_O[5]/FROM )
    );
    X_BUF \SDAT_O<5>/YUSED (
      .I (\SDAT_O[5]/GROM ),
      .O (syn178395)
    );
    X_BUF \SDAT_O<5>/XUSED (
      .I (\SDAT_O[5]/FROM ),
      .O (SDAT_O[5])
    );
    defparam C19543.INIT = 16'hF888;
    X_LUT4 C19543(
      .ADR0 (\bridge/configuration/pci_err_addr [5]),
      .ADR1 (syn16984),
      .ADR2 (syn17074),
      .ADR3 (\bridge/configuration/wb_err_data [5]),
      .O (\syn178393/GROM )
    );
    defparam C19542.INIT = 16'hF8F8;
    X_LUT4 C19542(
      .ADR0 (syn17084),
      .ADR1 (\bridge/configuration/interrupt_line [5]),
      .ADR2 (syn178390),
      .ADR3 (VCC),
      .O (\syn178393/FROM )
    );
    X_BUF \syn178393/YUSED (
      .I (\syn178393/GROM ),
      .O (syn178390)
    );
    X_BUF \syn178393/XUSED (
      .I (\syn178393/FROM ),
      .O (syn178393)
    );
    defparam C19586.INIT = 16'hAA00;
    X_LUT4 C19586(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn178392/GROM )
    );
    defparam C19540.INIT = 16'hF888;
    X_LUT4 C19540(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [5]),
      .ADR1 (syn17745),
      .ADR2 (syn17078),
      .ADR3 (\bridge/configuration/wb_err_addr [5]),
      .O (\syn178392/FROM )
    );
    X_BUF \syn178392/YUSED (
      .I (\syn178392/GROM ),
      .O (syn17078)
    );
    X_BUF \syn178392/XUSED (
      .I (\syn178392/FROM ),
      .O (syn178392)
    );
    defparam C19532.INIT = 16'hECA0;
    X_LUT4 C19532(
      .ADR0 (syn17083),
      .ADR1 (\bridge/configuration/pci_err_data [4]),
      .ADR2 (\bridge/configuration/interrupt_line [4]),
      .ADR3 (syn17072),
      .O (\SDAT_O[4]/GROM )
    );
    defparam C19531.INIT = 16'hFFFE;
    X_LUT4 C19531(
      .ADR0 (syn18717),
      .ADR1 (syn178410),
      .ADR2 (syn178411),
      .ADR3 (syn178409),
      .O (\SDAT_O[4]/FROM )
    );
    X_BUF \SDAT_O<4>/YUSED (
      .I (\SDAT_O[4]/GROM ),
      .O (syn178411)
    );
    X_BUF \SDAT_O<4>/XUSED (
      .I (\SDAT_O[4]/FROM ),
      .O (SDAT_O[4])
    );
    defparam C19534.INIT = 16'h8080;
    X_LUT4 C19534(
      .ADR0 (syn16917),
      .ADR1 (\bridge/configuration/pci_err_addr [4]),
      .ADR2 (\bridge/configuration/C2338 ),
      .ADR3 (VCC),
      .O (\syn178410/GROM )
    );
    defparam C19533.INIT = 16'hFFF8;
    X_LUT4 C19533(
      .ADR0 (syn17745),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [4]),
      .ADR2 (syn18716),
      .ADR3 (syn18713),
      .O (\syn178410/FROM )
    );
    X_BUF \syn178410/YUSED (
      .I (\syn178410/GROM ),
      .O (syn18716)
    );
    X_BUF \syn178410/XUSED (
      .I (\syn178410/FROM ),
      .O (syn178410)
    );
    defparam C19522.INIT = 16'hFEFA;
    X_LUT4 C19522(
      .ADR0 (syn178432),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [3]),
      .ADR2 (syn178433),
      .ADR3 (syn17745),
      .O (\SDAT_O[3]/GROM )
    );
    defparam C19521.INIT = 16'hAAA8;
    X_LUT4 C19521(
      .ADR0 (syn24476),
      .ADR1 (syn178436),
      .ADR2 (syn178437),
      .ADR3 (syn178435),
      .O (\SDAT_O[3]/FROM )
    );
    X_BUF \SDAT_O<3>/YUSED (
      .I (\SDAT_O[3]/GROM ),
      .O (syn178437)
    );
    X_BUF \SDAT_O<3>/XUSED (
      .I (\SDAT_O[3]/FROM ),
      .O (SDAT_O[3])
    );
    defparam C19527.INIT = 16'h8000;
    X_LUT4 C19527(
      .ADR0 (syn177458),
      .ADR1 (syn177397),
      .ADR2 (\bridge/configuration/serr_int_en ),
      .ADR3 (syn177396),
      .O (\syn178435/GROM )
    );
    defparam C19526.INIT = 16'hEAC0;
    X_LUT4 C19526(
      .ADR0 (syn17084),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR2 (syn18725),
      .ADR3 (\bridge/configuration/interrupt_line [3]),
      .O (\syn178435/FROM )
    );
    X_BUF \syn178435/YUSED (
      .I (\syn178435/GROM ),
      .O (syn18725)
    );
    X_BUF \syn178435/XUSED (
      .I (\syn178435/FROM ),
      .O (syn178435)
    );
    defparam C19596.INIT = 16'hF000;
    X_LUT4 C19596(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR3 (\bridge/configuration/C2302 ),
      .O (\syn178432/GROM )
    );
    defparam C19524.INIT = 16'hF888;
    X_LUT4 C19524(
      .ADR0 (syn16984),
      .ADR1 (\bridge/configuration/pci_err_addr [3]),
      .ADR2 (syn17074),
      .ADR3 (\bridge/configuration/wb_err_data [3]),
      .O (\syn178432/FROM )
    );
    X_BUF \syn178432/YUSED (
      .I (\syn178432/GROM ),
      .O (syn17074)
    );
    X_BUF \syn178432/XUSED (
      .I (\syn178432/FROM ),
      .O (syn178432)
    );
    defparam C19510.INIT = 16'hEAC0;
    X_LUT4 C19510(
      .ADR0 (\bridge/configuration/interrupt_line [2]),
      .ADR1 (syn17067),
      .ADR2 (\bridge/conf_cache_line_size_out [2]),
      .ADR3 (syn17083),
      .O (\SDAT_O[2]/GROM )
    );
    defparam C19509.INIT = 16'hFEFA;
    X_LUT4 C19509(
      .ADR0 (syn178469),
      .ADR1 (syn16917),
      .ADR2 (syn178470),
      .ADR3 (syn18765),
      .O (\SDAT_O[2]/FROM )
    );
    X_BUF \SDAT_O<2>/YUSED (
      .I (\SDAT_O[2]/GROM ),
      .O (syn178470)
    );
    X_BUF \SDAT_O<2>/XUSED (
      .I (\SDAT_O[2]/FROM ),
      .O (SDAT_O[2])
    );
    defparam C19513.INIT = 16'hFEFE;
    X_LUT4 C19513(
      .ADR0 (syn178459),
      .ADR1 (syn178462),
      .ADR2 (syn178460),
      .ADR3 (VCC),
      .O (\syn18765/GROM )
    );
    defparam C19512.INIT = 16'hFFF8;
    X_LUT4 C19512(
      .ADR0 (\bridge/configuration/C2334 ),
      .ADR1 (\bridge/configuration/pci_err_data [2]),
      .ADR2 (syn178465),
      .ADR3 (syn18756),
      .O (\syn18765/FROM )
    );
    X_BUF \syn18765/YUSED (
      .I (\syn18765/GROM ),
      .O (syn178465)
    );
    X_BUF \syn18765/XUSED (
      .I (\syn18765/FROM ),
      .O (syn18765)
    );
    defparam C19517.INIT = 16'h8080;
    X_LUT4 C19517(
      .ADR0 (syn178449),
      .ADR1 (syn177397),
      .ADR2 (syn177396),
      .ADR3 (VCC),
      .O (\syn178459/GROM )
    );
    defparam C19516.INIT = 16'hF888;
    X_LUT4 C19516(
      .ADR0 (\bridge/configuration/perr_int_en ),
      .ADR1 (\bridge/configuration/C2292 ),
      .ADR2 (\bridge/configuration/C2326 ),
      .ADR3 (\bridge/configuration/wb_img_ctrl1[2] ),
      .O (\syn178459/FROM )
    );
    X_BUF \syn178459/YUSED (
      .I (\syn178459/GROM ),
      .O (\bridge/configuration/C2326 )
    );
    X_BUF \syn178459/XUSED (
      .I (\syn178459/FROM ),
      .O (syn178459)
    );
    defparam C19927.INIT = 16'h0033;
    X_LUT4 C19927(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .O (\syn178449/GROM )
    );
    defparam C19518.INIT = 16'h2000;
    X_LUT4 C19518(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR2 (syn177450),
      .ADR3 (syn60060),
      .O (\syn178449/FROM )
    );
    X_BUF \syn178449/YUSED (
      .I (\syn178449/GROM ),
      .O (syn177450)
    );
    X_BUF \syn178449/XUSED (
      .I (\syn178449/FROM ),
      .O (syn178449)
    );
    defparam C19502.INIT = 16'hCCC8;
    X_LUT4 C19502(
      .ADR0 (syn178488),
      .ADR1 (syn16917),
      .ADR2 (syn18784),
      .ADR3 (syn178489),
      .O (\SDAT_O[1]/GROM )
    );
    defparam C19499.INIT = 16'hFFFC;
    X_LUT4 C19499(
      .ADR0 (VCC),
      .ADR1 (syn178495),
      .ADR2 (syn18800),
      .ADR3 (syn178494),
      .O (\SDAT_O[1]/FROM )
    );
    X_BUF \SDAT_O<1>/YUSED (
      .I (\SDAT_O[1]/GROM ),
      .O (syn18800)
    );
    X_BUF \SDAT_O<1>/XUSED (
      .I (\SDAT_O[1]/FROM ),
      .O (SDAT_O[1])
    );
    defparam C19506.INIT = 16'hEAC0;
    X_LUT4 C19506(
      .ADR0 (\bridge/configuration/C2326 ),
      .ADR1 (\bridge/configuration/C2292 ),
      .ADR2 (\bridge/configuration/error_int_en ),
      .ADR3 (\bridge/conf_wb_img_ctrl1_out [1]),
      .O (\syn178488/GROM )
    );
    defparam C19505.INIT = 16'hFCF0;
    X_LUT4 C19505(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/wb_err_addr [1]),
      .ADR2 (syn178485),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn178488/FROM )
    );
    X_BUF \syn178488/YUSED (
      .I (\syn178488/GROM ),
      .O (syn178485)
    );
    X_BUF \syn178488/XUSED (
      .I (\syn178488/FROM ),
      .O (syn178488)
    );
    defparam C19504.INIT = 16'hECA0;
    X_LUT4 C19504(
      .ADR0 (\bridge/configuration/wb_err_data [1]),
      .ADR1 (\bridge/configuration/C2338 ),
      .ADR2 (\bridge/configuration/C2302 ),
      .ADR3 (\bridge/configuration/pci_err_addr [1]),
      .O (\syn178489/GROM )
    );
    defparam C19503.INIT = 16'hF8F8;
    X_LUT4 C19503(
      .ADR0 (\bridge/configuration/pci_err_data [1]),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (syn178486),
      .ADR3 (VCC),
      .O (\syn178489/FROM )
    );
    X_BUF \syn178489/YUSED (
      .I (\syn178489/GROM ),
      .O (syn178486)
    );
    X_BUF \syn178489/XUSED (
      .I (\syn178489/FROM ),
      .O (syn178489)
    );
    defparam C19487.INIT = 16'hFFFA;
    X_LUT4 C19487(
      .ADR0 (syn178530),
      .ADR1 (VCC),
      .ADR2 (syn178529),
      .ADR3 (syn178528),
      .O (\SDAT_O[0]/GROM )
    );
    defparam C19486.INIT = 16'hFAF8;
    X_LUT4 C19486(
      .ADR0 (syn16917),
      .ADR1 (syn178523),
      .ADR2 (syn178532),
      .ADR3 (syn178522),
      .O (\SDAT_O[0]/FROM )
    );
    X_BUF \SDAT_O<0>/YUSED (
      .I (\SDAT_O[0]/GROM ),
      .O (syn178532)
    );
    X_BUF \SDAT_O<0>/XUSED (
      .I (\SDAT_O[0]/FROM ),
      .O (SDAT_O[0])
    );
    defparam C19492.INIT = 16'hFCCC;
    X_LUT4 C19492(
      .ADR0 (VCC),
      .ADR1 (syn178516),
      .ADR2 (\bridge/configuration/pci_err_data [0]),
      .ADR3 (\bridge/configuration/C2334 ),
      .O (\syn178523/GROM )
    );
    defparam C19491.INIT = 16'hFEFA;
    X_LUT4 C19491(
      .ADR0 (syn178517),
      .ADR1 (\bridge/configuration/pci_error_en ),
      .ADR2 (syn178520),
      .ADR3 (\bridge/configuration/C2340 ),
      .O (\syn178523/FROM )
    );
    X_BUF \syn178523/YUSED (
      .I (\syn178523/GROM ),
      .O (syn178520)
    );
    X_BUF \syn178523/XUSED (
      .I (\syn178523/FROM ),
      .O (syn178523)
    );
    defparam C19445.INIT = 16'h4400;
    X_LUT4 C19445(
      .ADR0 (syn17008),
      .ADR1 (syn18944),
      .ADR2 (VCC),
      .ADR3 (N12607),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N35/GROM )
    );
    defparam C19444.INIT = 16'hEAC0;
    X_LUT4 C19444(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [5])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [5]),
      .ADR2 (syn17085),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N35/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N35/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N35/GROM ),
      .O (syn17085)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N35/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N35/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N35 )
    );
    defparam C19977.INIT = 16'h8000;
    X_LUT4 C19977(
      .ADR0 (syn17678),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/C707 ),
      .ADR2 (syn177324),
      .ADR3 (\CRT/ssvga_wbm_if/S_41/cell0 ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow/GROM )
    );
    defparam C19447.INIT = 16'hF0F4;
    X_LUT4 C19447(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty ),
      .ADR1 (syn16935),
      .ADR2 (syn17008),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow/GROM ),
      .O (syn17008)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow )
    );
    defparam C19981.INIT = 16'h0008;
    X_LUT4 C19981(
      .ADR0 (syn177406),
      .ADR1 (syn177324),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/map ),
      .ADR3 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .O (\syn16935/GROM )
    );
    defparam C19980.INIT = 16'h8000;
    X_LUT4 C19980(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/img_hit [0]),
      .ADR1 (syn17669),
      .ADR2 (syn177343),
      .ADR3 (\CRT/ssvga_wbm_if/S_41/cell0 ),
      .O (\syn16935/FROM )
    );
    X_BUF \syn16935/YUSED (
      .I (\syn16935/GROM ),
      .O (syn177343)
    );
    X_BUF \syn16935/XUSED (
      .I (\syn16935/FROM ),
      .O (syn16935)
    );
    defparam C19990.INIT = 16'hFEFE;
    X_LUT4 C19990(
      .ADR0 (syn176894),
      .ADR1 (syn176895),
      .ADR2 (syn177317),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/S_41/cell0/GROM )
    );
    defparam C19988.INIT = 16'hAAA8;
    X_LUT4 C19988(
      .ADR0 (syn177324),
      .ADR1 (syn177319),
      .ADR2 (syn177321),
      .ADR3 (syn177320),
      .O (\CRT/ssvga_wbm_if/S_41/cell0/FROM )
    );
    X_BUF \CRT/ssvga_wbm_if/S_41/cell0/YUSED (
      .I (\CRT/ssvga_wbm_if/S_41/cell0/GROM ),
      .O (syn177321)
    );
    X_BUF \CRT/ssvga_wbm_if/S_41/cell0/XUSED (
      .I (\CRT/ssvga_wbm_if/S_41/cell0/FROM ),
      .O (\CRT/ssvga_wbm_if/S_41/cell0 )
    );
    defparam C19997.INIT = 16'h0FF0;
    X_LUT4 C19997(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [2]),
      .ADR3 (\CRT/ssvga_fifo/gray_read_ptr [4]),
      .O (\syn177319/GROM )
    );
    defparam C19996.INIT = 16'hDB7E;
    X_LUT4 C19996(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr_plus1 [3]),
      .ADR1 (\CRT/ssvga_fifo/gray_read_ptr [5]),
      .ADR2 (syn177311),
      .ADR3 (\CRT/ssvga_fifo/wr_ptr_plus1 [4]),
      .O (\syn177319/FROM )
    );
    X_BUF \syn177319/YUSED (
      .I (\syn177319/GROM ),
      .O (syn177311)
    );
    X_BUF \syn177319/XUSED (
      .I (\syn177319/FROM ),
      .O (syn177319)
    );
    defparam C19995.INIT = 16'h5A5A;
    X_LUT4 C19995(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr_plus1 [0]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/gray_read_ptr [2]),
      .ADR3 (VCC),
      .O (\syn177320/GROM )
    );
    defparam C19994.INIT = 16'hBD7E;
    X_LUT4 C19994(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr_plus1 [2]),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [1]),
      .ADR2 (syn177315),
      .ADR3 (\CRT/ssvga_fifo/gray_read_ptr [3]),
      .O (\syn177320/FROM )
    );
    X_BUF \syn177320/YUSED (
      .I (\syn177320/GROM ),
      .O (syn177315)
    );
    X_BUF \syn177320/XUSED (
      .I (\syn177320/FROM ),
      .O (syn177320)
    );
    defparam C19442.INIT = 16'h0100;
    X_LUT4 C19442(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_full_out ),
      .ADR1 (syn177324),
      .ADR2 (N12360),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [4]),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N30/GROM )
    );
    defparam C19441.INIT = 16'hFEFA;
    X_LUT4 C19441(
      .ADR0 (syn18958),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [4]),
      .ADR2 (syn18959),
      .ADR3 (syn17085),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N30/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N30/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N30/GROM ),
      .O (syn18959)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N30/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N30/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N30 )
    );
    defparam C19439.INIT = 16'h3300;
    X_LUT4 C19439(
      .ADR0 (VCC),
      .ADR1 (N12607),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [3]),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N24/GROM )
    );
    defparam C19438.INIT = 16'hFEFA;
    X_LUT4 C19438(
      .ADR0 (syn18965),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [3]),
      .ADR2 (syn18966),
      .ADR3 (syn17085),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N24/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N24/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N24/GROM ),
      .O (syn18966)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N24/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N24/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N24 )
    );
    defparam C19436.INIT = 16'h3030;
    X_LUT4 C19436(
      .ADR0 (VCC),
      .ADR1 (N12607),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [2]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N18/GROM )
    );
    defparam C19435.INIT = 16'hFFF8;
    X_LUT4 C19435(
      .ADR0 (syn17085),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [2]),
      .ADR2 (syn18973),
      .ADR3 (syn18972),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N18/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N18/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N18/GROM ),
      .O (syn18973)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N18/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N18/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N18 )
    );
    defparam C19433.INIT = 16'h5050;
    X_LUT4 C19433(
      .ADR0 (N12607),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [1]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N12/GROM )
    );
    defparam C19432.INIT = 16'hFEFA;
    X_LUT4 C19432(
      .ADR0 (syn18979),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [1]),
      .ADR2 (syn18980),
      .ADR3 (syn17085),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N12/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N12/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N12/GROM ),
      .O (syn18980)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N12/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N12/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N12 )
    );
    defparam C19430.INIT = 16'h5500;
    X_LUT4 C19430(
      .ADR0 (N12607),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_waddr [0]),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N6/GROM )
    );
    defparam C19429.INIT = 16'hFEFA;
    X_LUT4 C19429(
      .ADR0 (syn18984),
      .ADR1 (syn17085),
      .ADR2 (syn18985),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [0]),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N6/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N6/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N6/GROM ),
      .O (syn18985)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C6/N6/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C6/N6/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C6/N6 )
    );
    defparam C19299.INIT = 16'hFF80;
    X_LUT4 C19299(
      .ADR0 (syn17000),
      .ADR1 (syn24519),
      .ADR2 (syn24524),
      .ADR3 (syn178898),
      .O (\bridge/pci_target_unit/fifos/pcir_rallow/GROM )
    );
    defparam C19298.INIT = 16'hF000;
    X_LUT4 C19298(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn19420),
      .ADR3 (syn19407),
      .O (\bridge/pci_target_unit/fifos/pcir_rallow/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_rallow/YUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_rallow/GROM ),
      .O (syn19420)
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_rallow/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_rallow/FROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_rallow )
    );
    defparam C19294.INIT = 16'h0CAA;
    X_LUT4 C19294(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_waddr [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_raddr [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR3 (N12616),
      .O (\bridge/pci_target_unit/fifos/C9/N30/GROM )
    );
    defparam C19293.INIT = 16'hF8F0;
    X_LUT4 C19293(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_raddr_0 [4]),
      .ADR2 (syn178911),
      .ADR3 (N12616),
      .O (\bridge/pci_target_unit/fifos/C9/N30/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N30/YUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N30/GROM ),
      .O (syn178911)
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N30/XUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N30/FROM ),
      .O (\bridge/pci_target_unit/fifos/C9/N30 )
    );
    defparam C19291.INIT = 16'h0CAC;
    X_LUT4 C19291(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_raddr [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_waddr [3]),
      .ADR2 (N12616),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .O (\bridge/pci_target_unit/fifos/C9/N24/GROM )
    );
    defparam C19290.INIT = 16'hF8F0;
    X_LUT4 C19290(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_raddr_0 [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR2 (syn178919),
      .ADR3 (N12616),
      .O (\bridge/pci_target_unit/fifos/C9/N24/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N24/YUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N24/GROM ),
      .O (syn178919)
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N24/XUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N24/FROM ),
      .O (\bridge/pci_target_unit/fifos/C9/N24 )
    );
    defparam C19288.INIT = 16'h4E44;
    X_LUT4 C19288(
      .ADR0 (N12616),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_waddr [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_raddr [2]),
      .O (\bridge/pci_target_unit/fifos/C9/N18/GROM )
    );
    defparam C19287.INIT = 16'hF8F0;
    X_LUT4 C19287(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_raddr_0 [2]),
      .ADR2 (syn178927),
      .ADR3 (N12616),
      .O (\bridge/pci_target_unit/fifos/C9/N18/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N18/YUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N18/GROM ),
      .O (syn178927)
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N18/XUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N18/FROM ),
      .O (\bridge/pci_target_unit/fifos/C9/N18 )
    );
    defparam C19285.INIT = 16'h3B08;
    X_LUT4 C19285(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_raddr [1]),
      .ADR1 (N12616),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_waddr [1]),
      .O (\bridge/pci_target_unit/fifos/C9/N12/GROM )
    );
    defparam C19284.INIT = 16'hF8F0;
    X_LUT4 C19284(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR1 (N12616),
      .ADR2 (syn178935),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_raddr_0 [1]),
      .O (\bridge/pci_target_unit/fifos/C9/N12/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N12/YUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N12/GROM ),
      .O (syn178935)
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N12/XUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N12/FROM ),
      .O (\bridge/pci_target_unit/fifos/C9/N12 )
    );
    defparam C19282.INIT = 16'h2F20;
    X_LUT4 C19282(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_raddr [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR2 (N12616),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_waddr [0]),
      .O (\bridge/pci_target_unit/fifos/C9/N6/GROM )
    );
    defparam C19281.INIT = 16'hF8F0;
    X_LUT4 C19281(
      .ADR0 (N12616),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_write_performed ),
      .ADR2 (syn178943),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_raddr_0 [0]),
      .O (\bridge/pci_target_unit/fifos/C9/N6/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N6/YUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N6/GROM ),
      .O (syn178943)
    );
    X_BUF \bridge/pci_target_unit/fifos/C9/N6/XUSED (
      .I (\bridge/pci_target_unit/fifos/C9/N6/FROM ),
      .O (\bridge/pci_target_unit/fifos/C9/N6 )
    );
    defparam C19168.INIT = 16'hC3FF;
    X_LUT4 C19168(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_pci_ba1_out [15]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .ADR3 (\bridge/conf_pci_am1_out [15]),
      .O (\syn179246/GROM )
    );
    defparam C19167.INIT = 16'h90F0;
    X_LUT4 C19167(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .ADR1 (\bridge/conf_pci_ba1_out [16]),
      .ADR2 (syn19873),
      .ADR3 (\bridge/conf_pci_am1_out [16]),
      .O (\syn179246/FROM )
    );
    X_BUF \syn179246/YUSED (
      .I (\syn179246/GROM ),
      .O (syn19873)
    );
    X_BUF \syn179246/XUSED (
      .I (\syn179246/FROM ),
      .O (syn179246)
    );
    defparam C19166.INIT = 16'h9F9F;
    X_LUT4 C19166(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .ADR1 (\bridge/conf_pci_ba1_out [13]),
      .ADR2 (\bridge/conf_pci_am1_out [13]),
      .ADR3 (VCC),
      .O (\syn179247/GROM )
    );
    defparam C19165.INIT = 16'h90F0;
    X_LUT4 C19165(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .ADR1 (\bridge/conf_pci_ba1_out [14]),
      .ADR2 (syn19881),
      .ADR3 (\bridge/conf_pci_am1_out [14]),
      .O (\syn179247/FROM )
    );
    X_BUF \syn179247/YUSED (
      .I (\syn179247/GROM ),
      .O (syn19881)
    );
    X_BUF \syn179247/XUSED (
      .I (\syn179247/FROM ),
      .O (syn179247)
    );
    defparam C19164.INIT = 16'hF0CC;
    X_LUT4 C19164(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_mem_space_enable_out ),
      .ADR2 (\bridge/conf_io_space_enable_out ),
      .ADR3 (\bridge/conf_pci_mem_io1_out ),
      .O (\syn179248/GROM )
    );
    defparam C19163.INIT = 16'hD070;
    X_LUT4 C19163(
      .ADR0 (\bridge/conf_pci_am1_out [12]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .ADR2 (syn19884),
      .ADR3 (\bridge/conf_pci_ba1_out [12]),
      .O (\syn179248/FROM )
    );
    X_BUF \syn179248/YUSED (
      .I (\syn179248/GROM ),
      .O (syn19884)
    );
    X_BUF \syn179248/XUSED (
      .I (\syn179248/FROM ),
      .O (syn179248)
    );
    defparam C19142.INIT = 16'hCCD8;
    X_LUT4 C19142(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg [1]),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_control_out [1]),
      .ADR3 (\bridge/in_reg_irdy_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy/GROM )
    );
    defparam C19139.INIT = 16'hCC40;
    X_LUT4 C19139(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/N64 ),
      .ADR2 (\bridge/pci_target_unit/pcit_if_pcir_fifo_data_err_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_disconect_wo_data_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pcir_fifo_data_err_out )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy )
    );
    defparam C19145.INIT = 16'h0003;
    X_LUT4 C19145(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos_pciw_full_out ),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_full ),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_two_left_out ),
      .O (\syn179287/GROM )
    );
    defparam C19144.INIT = 16'hFFAE;
    X_LUT4 C19144(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/conf_addr_out [0]),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR2 (syn19927),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/conf_addr_out [1]),
      .O (\syn179287/FROM )
    );
    X_BUF \syn179287/YUSED (
      .I (\syn179287/GROM ),
      .O (syn19927)
    );
    X_BUF \syn179287/XUSED (
      .I (\syn179287/FROM ),
      .O (syn179287)
    );
    defparam C19133.INIT = 16'h0040;
    X_LUT4 C19133(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/N59 ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/same_read_reg ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/rd_progress ),
      .O (\syn19968/GROM )
    );
    defparam C19132.INIT = 16'h00F2;
    X_LUT4 C19132(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/wr_progress ),
      .ADR2 (syn19963),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/cnf_progress ),
      .O (\syn19968/FROM )
    );
    X_BUF \syn19968/YUSED (
      .I (\syn19968/GROM ),
      .O (syn19963)
    );
    X_BUF \syn19968/XUSED (
      .I (\syn19968/FROM ),
      .O (syn19968)
    );
    defparam C19975.INIT = 16'hAA22;
    X_LUT4 C19975(
      .ADR0 (\CRT/ssvga_wbm_if/S_41/cell0 ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_control_out [1]),
      .ADR2 (VCC),
      .ADR3 (syn17686),
      .O (\CRT/fifo_wr_en/GROM )
    );
    defparam C19974.INIT = 16'hF0E0;
    X_LUT4 C19974(
      .ADR0 (syn17686),
      .ADR1 (syn16935),
      .ADR2 (syn177358),
      .ADR3 (syn17008),
      .O (\CRT/fifo_wr_en/FROM )
    );
    X_BUF \CRT/fifo_wr_en/YUSED (
      .I (\CRT/fifo_wr_en/GROM ),
      .O (syn177358)
    );
    X_BUF \CRT/fifo_wr_en/XUSED (
      .I (\CRT/fifo_wr_en/FROM ),
      .O (\CRT/fifo_wr_en )
    );
    defparam C18772.INIT = 16'h2000;
    X_LUT4 C18772(
      .ADR0 (syn179659),
      .ADR1 (\bridge/pciu_conf_offset_out [2]),
      .ADR2 (syn60111),
      .ADR3 (\bridge/pciu_conf_offset_out [3]),
      .O (\syn17116/GROM )
    );
    defparam C18771.INIT = 16'hF000;
    X_LUT4 C18771(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/C2001 ),
      .ADR3 (syn16914),
      .O (\syn17116/FROM )
    );
    X_BUF \syn17116/YUSED (
      .I (\syn17116/GROM ),
      .O (\bridge/configuration/C2001 )
    );
    X_BUF \syn17116/XUSED (
      .I (\syn17116/FROM ),
      .O (syn17116)
    );
    defparam C19312.INIT = 16'h0505;
    X_LUT4 C19312(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/cnf_progress ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg ),
      .ADR3 (VCC),
      .O (\syn16914/GROM )
    );
    defparam C18780.INIT = 16'h0001;
    X_LUT4 C18780(
      .ADR0 (\bridge/out_bckp_devsel_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR2 (syn19366),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\syn16914/FROM )
    );
    X_BUF \syn16914/YUSED (
      .I (\syn16914/GROM ),
      .O (syn19366)
    );
    X_BUF \syn16914/XUSED (
      .I (\syn16914/FROM ),
      .O (syn16914)
    );
    defparam C18764.INIT = 16'hA000;
    X_LUT4 C18764(
      .ADR0 (syn17104),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/interrupt_line [0]),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn179881/GROM )
    );
    defparam C18763.INIT = 16'hF8F0;
    X_LUT4 C18763(
      .ADR0 (syn17101),
      .ADR1 (\bridge/conf_cache_line_size_out [0]),
      .ADR2 (syn20480),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn179881/FROM )
    );
    X_BUF \syn179881/YUSED (
      .I (\syn179881/GROM ),
      .O (syn20480)
    );
    X_BUF \syn179881/XUSED (
      .I (\syn179881/FROM ),
      .O (syn179881)
    );
    defparam C18694.INIT = 16'hFEEE;
    X_LUT4 C18694(
      .ADR0 (syn180051),
      .ADR1 (syn17121),
      .ADR2 (\bridge/configuration/interrupt_line [5]),
      .ADR3 (syn17105),
      .O (\syn20662/GROM )
    );
    defparam C18693.INIT = 16'hCCC8;
    X_LUT4 C18693(
      .ADR0 (syn180052),
      .ADR1 (syn180250),
      .ADR2 (syn180054),
      .ADR3 (syn180053),
      .O (\syn20662/FROM )
    );
    X_BUF \syn20662/YUSED (
      .I (\syn20662/GROM ),
      .O (syn180054)
    );
    X_BUF \syn20662/XUSED (
      .I (\syn20662/FROM ),
      .O (syn20662)
    );
    defparam C18728.INIT = 16'hF000;
    X_LUT4 C18728(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\syn180051/GROM )
    );
    defparam C18695.INIT = 16'hF888;
    X_LUT4 C18695(
      .ADR0 (\bridge/conf_cache_line_size_out [5]),
      .ADR1 (syn17102),
      .ADR2 (syn17016),
      .ADR3 (\bridge/configuration/config_addr[5] ),
      .O (\syn180051/FROM )
    );
    X_BUF \syn180051/YUSED (
      .I (\syn180051/GROM ),
      .O (syn17016)
    );
    X_BUF \syn180051/XUSED (
      .I (\syn180051/FROM ),
      .O (syn180051)
    );
    defparam C18905.INIT = 16'h5000;
    X_LUT4 C18905(
      .ADR0 (\bridge/pciu_conf_offset_out [4]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pciu_conf_offset_out [6]),
      .ADR3 (\bridge/pciu_conf_offset_out [5]),
      .O (\bridge/configuration/C1929/GROM )
    );
    defparam C18903.INIT = 16'h0020;
    X_LUT4 C18903(
      .ADR0 (\bridge/pciu_conf_offset_out [7]),
      .ADR1 (\bridge/pciu_conf_offset_out [2]),
      .ADR2 (syn17002),
      .ADR3 (\bridge/pciu_conf_offset_out [3]),
      .O (\bridge/configuration/C1929/FROM )
    );
    X_BUF \bridge/configuration/C1929/YUSED (
      .I (\bridge/configuration/C1929/GROM ),
      .O (syn17002)
    );
    X_BUF \bridge/configuration/C1929/XUSED (
      .I (\bridge/configuration/C1929/FROM ),
      .O (\bridge/configuration/C1929 )
    );
    defparam C18652.INIT = 16'h8000;
    X_LUT4 C18652(
      .ADR0 (syn60038),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn16985),
      .ADR3 (\bridge/configuration/pci_err_data [8]),
      .O (\syn180183/GROM )
    );
    defparam C18651.INIT = 16'hFFFE;
    X_LUT4 C18651(
      .ADR0 (syn20739),
      .ADR1 (syn20741),
      .ADR2 (syn20742),
      .ADR3 (syn20740),
      .O (\syn180183/FROM )
    );
    X_BUF \syn180183/YUSED (
      .I (\syn180183/GROM ),
      .O (syn20742)
    );
    X_BUF \syn180183/XUSED (
      .I (\syn180183/FROM ),
      .O (syn180183)
    );
    defparam C18664.INIT = 16'hFFAA;
    X_LUT4 C18664(
      .ADR0 (syn59991),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (syn17106),
      .O (\syn20739/GROM )
    );
    defparam C18655.INIT = 16'h8000;
    X_LUT4 C18655(
      .ADR0 (\bridge/configuration/config_addr[8] ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn60038),
      .ADR3 (syn17016),
      .O (\syn20739/FROM )
    );
    X_BUF \syn20739/YUSED (
      .I (\syn20739/GROM ),
      .O (syn60038)
    );
    X_BUF \syn20739/XUSED (
      .I (\syn20739/FROM ),
      .O (syn20739)
    );
    defparam C18794.INIT = 16'h8000;
    X_LUT4 C18794(
      .ADR0 (\bridge/pciu_conf_offset_out [6]),
      .ADR1 (syn17003),
      .ADR2 (\bridge/pciu_conf_offset_out [2]),
      .ADR3 (\bridge/pciu_conf_offset_out [7]),
      .O (\syn17015/GROM )
    );
    defparam C18729.INIT = 16'hF000;
    X_LUT4 C18729(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/C1935 ),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\syn17015/FROM )
    );
    X_BUF \syn17015/YUSED (
      .I (\syn17015/GROM ),
      .O (\bridge/configuration/C1935 )
    );
    X_BUF \syn17015/XUSED (
      .I (\syn17015/FROM ),
      .O (syn17015)
    );
    defparam C18792.INIT = 16'h0080;
    X_LUT4 C18792(
      .ADR0 (\bridge/pciu_conf_offset_out [6]),
      .ADR1 (syn17003),
      .ADR2 (\bridge/pciu_conf_offset_out [7]),
      .ADR3 (\bridge/pciu_conf_offset_out [2]),
      .O (\syn17014/GROM )
    );
    defparam C18725.INIT = 16'hC0C0;
    X_LUT4 C18725(
      .ADR0 (VCC),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1937 ),
      .ADR3 (VCC),
      .O (\syn17014/FROM )
    );
    X_BUF \syn17014/YUSED (
      .I (\syn17014/GROM ),
      .O (\bridge/configuration/C1937 )
    );
    X_BUF \syn17014/XUSED (
      .I (\syn17014/FROM ),
      .O (syn17014)
    );
    defparam C18798.INIT = 16'h0C00;
    X_LUT4 C18798(
      .ADR0 (VCC),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (\bridge/pciu_conf_offset_out [2]),
      .ADR3 (syn17103),
      .O (\syn16985/GROM )
    );
    defparam C18726.INIT = 16'hC0C0;
    X_LUT4 C18726(
      .ADR0 (VCC),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (VCC),
      .O (\syn16985/FROM )
    );
    X_BUF \syn16985/YUSED (
      .I (\syn16985/GROM ),
      .O (\bridge/configuration/C1967 )
    );
    X_BUF \syn16985/XUSED (
      .I (\syn16985/FROM ),
      .O (syn16985)
    );
    defparam C18882.INIT = 16'hC000;
    X_LUT4 C18882(
      .ADR0 (VCC),
      .ADR1 (syn60089),
      .ADR2 (\bridge/pciu_conf_offset_out [7]),
      .ADR3 (\bridge/pciu_conf_offset_out [6]),
      .O (\syn180247/GROM )
    );
    defparam C18628.INIT = 16'hFFEC;
    X_LUT4 C18628(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (syn180244),
      .ADR2 (\bridge/configuration/C1941 ),
      .ADR3 (syn20796),
      .O (\syn180247/FROM )
    );
    X_BUF \syn180247/YUSED (
      .I (\syn180247/GROM ),
      .O (\bridge/configuration/C1941 )
    );
    X_BUF \syn180247/XUSED (
      .I (\syn180247/FROM ),
      .O (syn180247)
    );
    defparam C18877.INIT = 16'h1010;
    X_LUT4 C18877(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (syn17103),
      .ADR3 (VCC),
      .O (\syn180240/GROM )
    );
    defparam C18629.INIT = 16'hECCC;
    X_LUT4 C18629(
      .ADR0 (\bridge/configuration/pci_error_rty_exp_set ),
      .ADR1 (syn180244),
      .ADR2 (\bridge/configuration/C1973 ),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\syn180240/FROM )
    );
    X_BUF \syn180240/YUSED (
      .I (\syn180240/GROM ),
      .O (\bridge/configuration/C1973 )
    );
    X_BUF \syn180240/XUSED (
      .I (\syn180240/FROM ),
      .O (syn180240)
    );
    defparam C18626.INIT = 16'hF888;
    X_LUT4 C18626(
      .ADR0 (syn17014),
      .ADR1 (\bridge/configuration/wb_err_addr [10]),
      .ADR2 (syn17015),
      .ADR3 (\bridge/configuration/wb_err_data [10]),
      .O (\syn180248/GROM )
    );
    defparam C18625.INIT = 16'hFEFA;
    X_LUT4 C18625(
      .ADR0 (syn20803),
      .ADR1 (\bridge/configuration/pci_err_data [10]),
      .ADR2 (syn180245),
      .ADR3 (syn16985),
      .O (\syn180248/FROM )
    );
    X_BUF \syn180248/YUSED (
      .I (\syn180248/GROM ),
      .O (syn180245)
    );
    X_BUF \syn180248/XUSED (
      .I (\syn180248/FROM ),
      .O (syn180248)
    );
    defparam C18563.INIT = 16'hFFFE;
    X_LUT4 C18563(
      .ADR0 (syn180418),
      .ADR1 (syn180417),
      .ADR2 (syn180419),
      .ADR3 (syn180420),
      .O (\syn20947/GROM )
    );
    defparam C18562.INIT = 16'hFFFE;
    X_LUT4 C18562(
      .ADR0 (syn48754),
      .ADR1 (syn20934),
      .ADR2 (syn180425),
      .ADR3 (syn180416),
      .O (\syn20947/FROM )
    );
    X_BUF \syn20947/YUSED (
      .I (\syn20947/GROM ),
      .O (syn180425)
    );
    X_BUF \syn20947/XUSED (
      .I (\syn20947/FROM ),
      .O (syn20947)
    );
    defparam C18870.INIT = 16'h0020;
    X_LUT4 C18870(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [6]),
      .ADR2 (syn17003),
      .ADR3 (\bridge/pciu_conf_offset_out [7]),
      .O (\syn180417/GROM )
    );
    defparam C18567.INIT = 16'hECA0;
    X_LUT4 C18567(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [14]),
      .ADR1 (\bridge/configuration/C1989 ),
      .ADR2 (\bridge/configuration/C1987 ),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [14]),
      .O (\syn180417/FROM )
    );
    X_BUF \syn180417/YUSED (
      .I (\syn180417/GROM ),
      .O (\bridge/configuration/C1987 )
    );
    X_BUF \syn180417/XUSED (
      .I (\syn180417/FROM ),
      .O (syn180417)
    );
    defparam C18872.INIT = 16'h3000;
    X_LUT4 C18872(
      .ADR0 (VCC),
      .ADR1 (\bridge/pciu_conf_offset_out [5]),
      .ADR2 (\bridge/pciu_conf_offset_out [4]),
      .ADR3 (\bridge/pciu_conf_offset_out [3]),
      .O (\bridge/configuration/C1989/GROM )
    );
    defparam C18871.INIT = 16'h0010;
    X_LUT4 C18871(
      .ADR0 (\bridge/pciu_conf_offset_out [6]),
      .ADR1 (\bridge/pciu_conf_offset_out [7]),
      .ADR2 (syn17003),
      .ADR3 (\bridge/pciu_conf_offset_out [2]),
      .O (\bridge/configuration/C1989/FROM )
    );
    X_BUF \bridge/configuration/C1989/YUSED (
      .I (\bridge/configuration/C1989/GROM ),
      .O (syn17003)
    );
    X_BUF \bridge/configuration/C1989/XUSED (
      .I (\bridge/configuration/C1989/FROM ),
      .O (\bridge/configuration/C1989 )
    );
    defparam C18910.INIT = 16'h0800;
    X_LUT4 C18910(
      .ADR0 (syn179659),
      .ADR1 (\bridge/pciu_conf_offset_out [2]),
      .ADR2 (\bridge/pciu_conf_offset_out [3]),
      .ADR3 (syn60111),
      .O (\syn180418/GROM )
    );
    defparam C18566.INIT = 16'hF888;
    X_LUT4 C18566(
      .ADR0 (\bridge/configuration/config_addr[14] ),
      .ADR1 (\bridge/configuration/C1929 ),
      .ADR2 (\bridge/configuration/C2003 ),
      .ADR3 (\bridge/configuration/pci_base_addr0 [14]),
      .O (\syn180418/FROM )
    );
    X_BUF \syn180418/YUSED (
      .I (\syn180418/GROM ),
      .O (\bridge/configuration/C2003 )
    );
    X_BUF \syn180418/XUSED (
      .I (\syn180418/FROM ),
      .O (syn180418)
    );
    defparam C18878.INIT = 16'h0200;
    X_LUT4 C18878(
      .ADR0 (\bridge/pciu_conf_offset_out [5]),
      .ADR1 (\bridge/pciu_conf_offset_out [7]),
      .ADR2 (\bridge/pciu_conf_offset_out [4]),
      .ADR3 (\bridge/pciu_conf_offset_out [6]),
      .O (\bridge/configuration/C1971/GROM )
    );
    defparam C18799.INIT = 16'h4040;
    X_LUT4 C18799(
      .ADR0 (\bridge/pciu_conf_offset_out [3]),
      .ADR1 (\bridge/pciu_conf_offset_out [2]),
      .ADR2 (syn17103),
      .ADR3 (VCC),
      .O (\bridge/configuration/C1971/FROM )
    );
    X_BUF \bridge/configuration/C1971/YUSED (
      .I (\bridge/configuration/C1971/GROM ),
      .O (syn17103)
    );
    X_BUF \bridge/configuration/C1971/XUSED (
      .I (\bridge/configuration/C1971/FROM ),
      .O (\bridge/configuration/C1971 )
    );
    defparam C18559.INIT = 16'hC000;
    X_LUT4 C18559(
      .ADR0 (VCC),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (\bridge/configuration/pci_base_addr0 [14]),
      .ADR3 (syn16929),
      .O (\syn180440/GROM )
    );
    defparam C18558.INIT = 16'hF8F0;
    X_LUT4 C18558(
      .ADR0 (syn17101),
      .ADR1 (\bridge/conf_latency_tim_out [6]),
      .ADR2 (syn20953),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn180440/FROM )
    );
    X_BUF \syn180440/YUSED (
      .I (\syn180440/GROM ),
      .O (syn20953)
    );
    X_BUF \syn180440/XUSED (
      .I (\syn180440/FROM ),
      .O (syn180440)
    );
    defparam C18884.INIT = 16'h0002;
    X_LUT4 C18884(
      .ADR0 (\bridge/pciu_conf_offset_out [4]),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (\bridge/pciu_conf_offset_out [5]),
      .ADR3 (\bridge/pciu_conf_offset_out [2]),
      .O (\syn16929/GROM )
    );
    defparam C18595.INIT = 16'h1000;
    X_LUT4 C18595(
      .ADR0 (\bridge/pciu_conf_offset_out [7]),
      .ADR1 (\bridge/pciu_conf_offset_out [6]),
      .ADR2 (syn60090),
      .ADR3 (syn16914),
      .O (\syn16929/FROM )
    );
    X_BUF \syn16929/YUSED (
      .I (\syn16929/GROM ),
      .O (syn60090)
    );
    X_BUF \syn16929/XUSED (
      .I (\syn16929/FROM ),
      .O (syn16929)
    );
    defparam C18546.INIT = 16'hFFFE;
    X_LUT4 C18546(
      .ADR0 (syn180470),
      .ADR1 (syn180469),
      .ADR2 (syn180468),
      .ADR3 (syn180467),
      .O (\syn20987/GROM )
    );
    defparam C18545.INIT = 16'hFFFE;
    X_LUT4 C18545(
      .ADR0 (syn20974),
      .ADR1 (syn48754),
      .ADR2 (syn180475),
      .ADR3 (syn180466),
      .O (\syn20987/FROM )
    );
    X_BUF \syn20987/YUSED (
      .I (\syn20987/GROM ),
      .O (syn180475)
    );
    X_BUF \syn20987/XUSED (
      .I (\syn20987/FROM ),
      .O (syn20987)
    );
    defparam C18542.INIT = 16'hA000;
    X_LUT4 C18542(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (VCC),
      .ADR2 (syn16929),
      .ADR3 (\bridge/configuration/pci_base_addr0 [15]),
      .O (\syn180490/GROM )
    );
    defparam C18541.INIT = 16'hF8F0;
    X_LUT4 C18541(
      .ADR0 (\bridge/conf_latency_tim_out [7]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn20993),
      .ADR3 (syn17101),
      .O (\syn180490/FROM )
    );
    X_BUF \syn180490/YUSED (
      .I (\syn180490/GROM ),
      .O (syn20993)
    );
    X_BUF \syn180490/XUSED (
      .I (\syn180490/FROM ),
      .O (syn180490)
    );
    defparam C18528.INIT = 16'hECA0;
    X_LUT4 C18528(
      .ADR0 (syn16929),
      .ADR1 (syn17065),
      .ADR2 (\bridge/configuration/pci_base_addr0 [16]),
      .ADR3 (syn16927),
      .O (\syn180535/GROM )
    );
    defparam C18527.INIT = 16'hFFFC;
    X_LUT4 C18527(
      .ADR0 (VCC),
      .ADR1 (syn17120),
      .ADR2 (syn180534),
      .ADR3 (syn180532),
      .O (\syn180535/FROM )
    );
    X_BUF \syn180535/YUSED (
      .I (\syn180535/GROM ),
      .O (syn180534)
    );
    X_BUF \syn180535/XUSED (
      .I (\syn180535/FROM ),
      .O (syn180535)
    );
    defparam C18915.INIT = 16'h0022;
    X_LUT4 C18915(
      .ADR0 (syn60089),
      .ADR1 (\bridge/pciu_conf_offset_out [7]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pciu_conf_offset_out [6]),
      .O (\syn16927/GROM )
    );
    defparam C18775.INIT = 16'h2020;
    X_LUT4 C18775(
      .ADR0 (syn17106),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (syn60110),
      .ADR3 (VCC),
      .O (\syn16927/FROM )
    );
    X_BUF \syn16927/YUSED (
      .I (\syn16927/GROM ),
      .O (syn60110)
    );
    X_BUF \syn16927/XUSED (
      .I (\syn16927/FROM ),
      .O (syn16927)
    );
    defparam C18510.INIT = 16'hECCC;
    X_LUT4 C18510(
      .ADR0 (syn17064),
      .ADR1 (syn180580),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn16927),
      .O (\syn180582/GROM )
    );
    defparam C18509.INIT = 16'hF8F0;
    X_LUT4 C18509(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn16929),
      .ADR2 (syn180581),
      .ADR3 (\bridge/configuration/pci_base_addr0 [17]),
      .O (\syn180582/FROM )
    );
    X_BUF \syn180582/YUSED (
      .I (\syn180582/GROM ),
      .O (syn180581)
    );
    X_BUF \syn180582/XUSED (
      .I (\syn180582/FROM ),
      .O (syn180582)
    );
    defparam C18768.INIT = 16'hA0A0;
    X_LUT4 C18768(
      .ADR0 (syn16919),
      .ADR1 (VCC),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (VCC),
      .O (\syn180580/GROM )
    );
    defparam C18511.INIT = 16'hF888;
    X_LUT4 C18511(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [17]),
      .ADR1 (syn136384),
      .ADR2 (syn136386),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [17]),
      .O (\syn180580/FROM )
    );
    X_BUF \syn180580/YUSED (
      .I (\syn180580/GROM ),
      .O (syn136386)
    );
    X_BUF \syn180580/XUSED (
      .I (\syn180580/FROM ),
      .O (syn180580)
    );
    defparam C18770.INIT = 16'h0032;
    X_LUT4 C18770(
      .ADR0 (\bridge/in_reg_irdy_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg ),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/cnf_progress ),
      .O (\syn136384/GROM )
    );
    defparam C18769.INIT = 16'hC0C0;
    X_LUT4 C18769(
      .ADR0 (VCC),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn16931),
      .ADR3 (VCC),
      .O (\syn136384/FROM )
    );
    X_BUF \syn136384/YUSED (
      .I (\syn136384/GROM ),
      .O (syn16931)
    );
    X_BUF \syn136384/XUSED (
      .I (\syn136384/FROM ),
      .O (syn136384)
    );
    defparam C18484.INIT = 16'hFFFE;
    X_LUT4 C18484(
      .ADR0 (syn180659),
      .ADR1 (syn180660),
      .ADR2 (syn180661),
      .ADR3 (syn180658),
      .O (\syn21143/GROM )
    );
    defparam C18483.INIT = 16'hFFFE;
    X_LUT4 C18483(
      .ADR0 (syn180657),
      .ADR1 (syn48754),
      .ADR2 (syn180666),
      .ADR3 (syn21130),
      .O (\syn21143/FROM )
    );
    X_BUF \syn21143/YUSED (
      .I (\syn21143/GROM ),
      .O (syn180666)
    );
    X_BUF \syn21143/XUSED (
      .I (\syn21143/FROM ),
      .O (syn21143)
    );
    defparam C18481.INIT = 16'hF888;
    X_LUT4 C18481(
      .ADR0 (syn16929),
      .ADR1 (\bridge/configuration/pci_base_addr0 [19]),
      .ADR2 (syn17062),
      .ADR3 (syn16927),
      .O (\syn180672/GROM )
    );
    defparam C18480.INIT = 16'hFFFA;
    X_LUT4 C18480(
      .ADR0 (syn180669),
      .ADR1 (VCC),
      .ADR2 (syn180671),
      .ADR3 (syn17104),
      .O (\syn180672/FROM )
    );
    X_BUF \syn180672/YUSED (
      .I (\syn180672/GROM ),
      .O (syn180671)
    );
    X_BUF \syn180672/XUSED (
      .I (\syn180672/FROM ),
      .O (syn180672)
    );
    defparam C18463.INIT = 16'hEAAA;
    X_LUT4 C18463(
      .ADR0 (syn180717),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn16927),
      .ADR3 (syn17061),
      .O (\syn180719/GROM )
    );
    defparam C18462.INIT = 16'hF8F0;
    X_LUT4 C18462(
      .ADR0 (\bridge/configuration/pci_base_addr0 [20]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180718),
      .ADR3 (syn16929),
      .O (\syn180719/FROM )
    );
    X_BUF \syn180719/YUSED (
      .I (\syn180719/GROM ),
      .O (syn180718)
    );
    X_BUF \syn180719/XUSED (
      .I (\syn180719/FROM ),
      .O (syn180719)
    );
    defparam C18447.INIT = 16'hECCC;
    X_LUT4 C18447(
      .ADR0 (syn16927),
      .ADR1 (syn180763),
      .ADR2 (syn17060),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn180765/GROM )
    );
    defparam C18446.INIT = 16'hF8F0;
    X_LUT4 C18446(
      .ADR0 (\bridge/configuration/pci_base_addr0 [21]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180764),
      .ADR3 (syn16929),
      .O (\syn180765/FROM )
    );
    X_BUF \syn180765/YUSED (
      .I (\syn180765/GROM ),
      .O (syn180764)
    );
    X_BUF \syn180765/XUSED (
      .I (\syn180765/FROM ),
      .O (syn180765)
    );
    defparam C18421.INIT = 16'hFFFE;
    X_LUT4 C18421(
      .ADR0 (syn180841),
      .ADR1 (syn180844),
      .ADR2 (syn180842),
      .ADR3 (syn180843),
      .O (\syn21298/GROM )
    );
    defparam C18420.INIT = 16'hFFFE;
    X_LUT4 C18420(
      .ADR0 (syn48754),
      .ADR1 (syn180840),
      .ADR2 (syn180849),
      .ADR3 (syn21285),
      .O (\syn21298/FROM )
    );
    X_BUF \syn21298/YUSED (
      .I (\syn21298/GROM ),
      .O (syn180849)
    );
    X_BUF \syn21298/XUSED (
      .I (\syn21298/FROM ),
      .O (syn21298)
    );
    defparam C18418.INIT = 16'hFEEE;
    X_LUT4 C18418(
      .ADR0 (syn17116),
      .ADR1 (syn180852),
      .ADR2 (syn16927),
      .ADR3 (syn17058),
      .O (\syn180855/GROM )
    );
    defparam C18417.INIT = 16'hF8F8;
    X_LUT4 C18417(
      .ADR0 (syn16929),
      .ADR1 (\bridge/configuration/pci_base_addr0 [23]),
      .ADR2 (syn180854),
      .ADR3 (VCC),
      .O (\syn180855/FROM )
    );
    X_BUF \syn180855/YUSED (
      .I (\syn180855/GROM ),
      .O (syn180854)
    );
    X_BUF \syn180855/XUSED (
      .I (\syn180855/FROM ),
      .O (syn180855)
    );
    defparam C18369.INIT = 16'hFFFE;
    X_LUT4 C18369(
      .ADR0 (syn181000),
      .ADR1 (syn180995),
      .ADR2 (syn180994),
      .ADR3 (syn181001),
      .O (\syn21430/GROM )
    );
    defparam C18365.INIT = 16'hEAEA;
    X_LUT4 C18365(
      .ADR0 (syn181008),
      .ADR1 (syn16916),
      .ADR2 (syn21421),
      .ADR3 (VCC),
      .O (\syn21430/FROM )
    );
    X_BUF \syn21430/YUSED (
      .I (\syn21430/GROM ),
      .O (syn21421)
    );
    X_BUF \syn21430/XUSED (
      .I (\syn21430/FROM ),
      .O (syn21430)
    );
    defparam C18375.INIT = 16'hECA0;
    X_LUT4 C18375(
      .ADR0 (\bridge/configuration/pci_err_addr [26]),
      .ADR1 (\bridge/configuration/pci_err_data [26]),
      .ADR2 (\bridge/configuration/C1971 ),
      .ADR3 (\bridge/configuration/C1967 ),
      .O (\syn181000/GROM )
    );
    defparam C18374.INIT = 16'hFFF8;
    X_LUT4 C18374(
      .ADR0 (\bridge/configuration/pci_err_cs_bit31_24 [26]),
      .ADR1 (\bridge/configuration/C1973 ),
      .ADR2 (syn180996),
      .ADR3 (syn48754),
      .O (\syn181000/FROM )
    );
    X_BUF \syn181000/YUSED (
      .I (\syn181000/GROM ),
      .O (syn180996)
    );
    X_BUF \syn181000/XUSED (
      .I (\syn181000/FROM ),
      .O (syn181000)
    );
    defparam C18371.INIT = 16'hECA0;
    X_LUT4 C18371(
      .ADR0 (\bridge/conf_pci_am1_out [14]),
      .ADR1 (\bridge/configuration/pci_tran_addr1 [26]),
      .ADR2 (\bridge/configuration/C1989 ),
      .ADR3 (\bridge/configuration/C1987 ),
      .O (\syn181001/GROM )
    );
    defparam C18370.INIT = 16'hFFFC;
    X_LUT4 C18370(
      .ADR0 (VCC),
      .ADR1 (syn180992),
      .ADR2 (syn180993),
      .ADR3 (syn21407),
      .O (\syn181001/FROM )
    );
    X_BUF \syn181001/YUSED (
      .I (\syn181001/GROM ),
      .O (syn180993)
    );
    X_BUF \syn181001/XUSED (
      .I (\syn181001/FROM ),
      .O (syn181001)
    );
    defparam C18900.INIT = 16'h4000;
    X_LUT4 C18900(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (syn179659),
      .ADR2 (\bridge/pciu_conf_offset_out [3]),
      .ADR3 (syn17004),
      .O (\syn21407/GROM )
    );
    defparam C18373.INIT = 16'hCC80;
    X_LUT4 C18373(
      .ADR0 (\bridge/conf_wb_ba1_out [14]),
      .ADR1 (\bridge/conf_wb_am1_out [14]),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/configuration/C1953 ),
      .O (\syn21407/FROM )
    );
    X_BUF \syn21407/YUSED (
      .I (\syn21407/GROM ),
      .O (\bridge/configuration/C1955 )
    );
    X_BUF \syn21407/XUSED (
      .I (\syn21407/FROM ),
      .O (syn21407)
    );
    defparam C18875.INIT = 16'h0008;
    X_LUT4 C18875(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (\bridge/pciu_conf_offset_out [4]),
      .ADR3 (\bridge/pciu_conf_offset_out [5]),
      .O (\bridge/configuration/C1953/GROM )
    );
    defparam C18874.INIT = 16'h2020;
    X_LUT4 C18874(
      .ADR0 (\bridge/pciu_conf_offset_out [7]),
      .ADR1 (\bridge/pciu_conf_offset_out [6]),
      .ADR2 (\bridge/configuration/C2268 ),
      .ADR3 (VCC),
      .O (\bridge/configuration/C1953/FROM )
    );
    X_BUF \bridge/configuration/C1953/YUSED (
      .I (\bridge/configuration/C1953/GROM ),
      .O (\bridge/configuration/C2268 )
    );
    X_BUF \bridge/configuration/C1953/XUSED (
      .I (\bridge/configuration/C1953/FROM ),
      .O (\bridge/configuration/C1953 )
    );
    defparam C18367.INIT = 16'hFEFC;
    X_LUT4 C18367(
      .ADR0 (syn17055),
      .ADR1 (syn181005),
      .ADR2 (syn17116),
      .ADR3 (syn16927),
      .O (\syn181008/GROM )
    );
    defparam C18366.INIT = 16'hFCF0;
    X_LUT4 C18366(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_pci_ba0_out [14]),
      .ADR2 (syn181007),
      .ADR3 (syn16929),
      .O (\syn181008/FROM )
    );
    X_BUF \syn181008/YUSED (
      .I (\syn181008/GROM ),
      .O (syn181007)
    );
    X_BUF \syn181008/XUSED (
      .I (\syn181008/FROM ),
      .O (syn181008)
    );
    defparam C18297.INIT = 16'hFEFE;
    X_LUT4 C18297(
      .ADR0 (syn181194),
      .ADR1 (syn181193),
      .ADR2 (syn21571),
      .ADR3 (VCC),
      .O (\syn21585/GROM )
    );
    defparam C18296.INIT = 16'hFFFE;
    X_LUT4 C18296(
      .ADR0 (syn181196),
      .ADR1 (syn181201),
      .ADR2 (syn181202),
      .ADR3 (syn181195),
      .O (\syn21585/FROM )
    );
    X_BUF \syn21585/YUSED (
      .I (\syn21585/GROM ),
      .O (syn181202)
    );
    X_BUF \syn21585/XUSED (
      .I (\syn21585/FROM ),
      .O (syn21585)
    );
    defparam C18302.INIT = 16'hEAC0;
    X_LUT4 C18302(
      .ADR0 (\bridge/configuration/pci_err_addr [30]),
      .ADR1 (\bridge/configuration/C1967 ),
      .ADR2 (\bridge/configuration/pci_err_data [30]),
      .ADR3 (\bridge/configuration/C1971 ),
      .O (\syn181201/GROM )
    );
    defparam C18301.INIT = 16'hFEFA;
    X_LUT4 C18301(
      .ADR0 (syn48754),
      .ADR1 (\bridge/configuration/C1973 ),
      .ADR2 (syn181197),
      .ADR3 (\bridge/configuration/pci_err_cs_bit31_24 [30]),
      .O (\syn181201/FROM )
    );
    X_BUF \syn181201/YUSED (
      .I (\syn181201/GROM ),
      .O (syn181197)
    );
    X_BUF \syn181201/XUSED (
      .I (\syn181201/FROM ),
      .O (syn181201)
    );
    defparam C18295.INIT = 16'h8000;
    X_LUT4 C18295(
      .ADR0 (syn16927),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (\bridge/conf_pci_am1_out [18]),
      .ADR3 (\bridge/conf_pci_ba1_out [18]),
      .O (\syn181217/GROM )
    );
    defparam C18294.INIT = 16'hF8F0;
    X_LUT4 C18294(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn17098),
      .ADR2 (syn21589),
      .ADR3 (\bridge/configuration/status_bit15_11 [14]),
      .O (\syn181217/FROM )
    );
    X_BUF \syn181217/YUSED (
      .I (\syn181217/GROM ),
      .O (syn21589)
    );
    X_BUF \syn181217/XUSED (
      .I (\syn181217/FROM ),
      .O (syn181217)
    );
    defparam C18278.INIT = 16'hFFFE;
    X_LUT4 C18278(
      .ADR0 (syn181251),
      .ADR1 (syn181250),
      .ADR2 (syn181249),
      .ADR3 (syn181252),
      .O (\syn21625/GROM )
    );
    defparam C18277.INIT = 16'hFFFE;
    X_LUT4 C18277(
      .ADR0 (syn181253),
      .ADR1 (syn181247),
      .ADR2 (syn181258),
      .ADR3 (syn181248),
      .O (\syn21625/FROM )
    );
    X_BUF \syn21625/YUSED (
      .I (\syn21625/GROM ),
      .O (syn181258)
    );
    X_BUF \syn21625/XUSED (
      .I (\syn21625/FROM ),
      .O (syn21625)
    );
    defparam C18276.INIT = 16'h8000;
    X_LUT4 C18276(
      .ADR0 (\bridge/conf_pci_ba1_out [19]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (\bridge/conf_pci_am1_out [19]),
      .ADR3 (syn16927),
      .O (\syn181272/GROM )
    );
    defparam C18275.INIT = 16'hF8F0;
    X_LUT4 C18275(
      .ADR0 (\bridge/configuration/status_bit15_11 [15]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn21629),
      .ADR3 (syn17098),
      .O (\syn181272/FROM )
    );
    X_BUF \syn181272/YUSED (
      .I (\syn181272/GROM ),
      .O (syn21629)
    );
    X_BUF \syn181272/XUSED (
      .I (\syn181272/FROM ),
      .O (syn181272)
    );
    defparam C18169.INIT = 16'h8222;
    X_LUT4 C18169(
      .ADR0 (syn181497),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [2]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR3 (syn24500),
      .O (\syn181520/GROM )
    );
    defparam C18168.INIT = 16'hC000;
    X_LUT4 C18168(
      .ADR0 (VCC),
      .ADR1 (syn181498),
      .ADR2 (syn181512),
      .ADR3 (syn181499),
      .O (\syn181520/FROM )
    );
    X_BUF \syn181520/YUSED (
      .I (\syn181520/GROM ),
      .O (syn181512)
    );
    X_BUF \syn181520/XUSED (
      .I (\syn181520/FROM ),
      .O (syn181520)
    );
    defparam C18176.INIT = 16'hC30F;
    X_LUT4 C18176(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [31]),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [31]),
      .ADR3 (syn24500),
      .O (\syn181498/GROM )
    );
    defparam C18175.INIT = 16'h8070;
    X_LUT4 C18175(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [29]),
      .ADR1 (syn24500),
      .ADR2 (syn176956),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [29]),
      .O (\syn181498/FROM )
    );
    X_BUF \syn181498/YUSED (
      .I (\syn181498/GROM ),
      .O (syn176956)
    );
    X_BUF \syn181498/XUSED (
      .I (\syn181498/FROM ),
      .O (syn181498)
    );
    defparam C18174.INIT = 16'hC333;
    X_LUT4 C18174(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [28]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [28]),
      .ADR3 (syn24500),
      .O (\syn181499/GROM )
    );
    defparam C18173.INIT = 16'h9030;
    X_LUT4 C18173(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [27]),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [27]),
      .ADR2 (syn176958),
      .ADR3 (syn24500),
      .O (\syn181499/FROM )
    );
    X_BUF \syn181499/YUSED (
      .I (\syn181499/GROM ),
      .O (syn176958)
    );
    X_BUF \syn181499/XUSED (
      .I (\syn181499/FROM ),
      .O (syn181499)
    );
    defparam C18172.INIT = 16'h8000;
    X_LUT4 C18172(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [2]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [1]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [3]),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [0]),
      .O (\syn181497/GROM )
    );
    defparam C18170.INIT = 16'h8070;
    X_LUT4 C18170(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [30]),
      .ADR1 (syn24500),
      .ADR2 (syn181495),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [30]),
      .O (\syn181497/FROM )
    );
    X_BUF \syn181497/YUSED (
      .I (\syn181497/GROM ),
      .O (syn181495)
    );
    X_BUF \syn181497/XUSED (
      .I (\syn181497/FROM ),
      .O (syn181497)
    );
    defparam C18160.INIT = 16'h820A;
    X_LUT4 C18160(
      .ADR0 (syn176967),
      .ADR1 (syn24500),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [20]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [20]),
      .O (\syn181521/GROM )
    );
    defparam C18159.INIT = 16'h8000;
    X_LUT4 C18159(
      .ADR0 (syn181501),
      .ADR1 (syn181502),
      .ADR2 (syn181503),
      .ADR3 (syn181500),
      .O (\syn181521/FROM )
    );
    X_BUF \syn181521/YUSED (
      .I (\syn181521/GROM ),
      .O (syn181503)
    );
    X_BUF \syn181521/XUSED (
      .I (\syn181521/FROM ),
      .O (syn181521)
    );
    defparam C18167.INIT = 16'h9393;
    X_LUT4 C18167(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [26]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [26]),
      .ADR3 (VCC),
      .O (\syn181500/GROM )
    );
    defparam C18166.INIT = 16'h9050;
    X_LUT4 C18166(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [25]),
      .ADR1 (syn24500),
      .ADR2 (syn176960),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [25]),
      .O (\syn181500/FROM )
    );
    X_BUF \syn181500/YUSED (
      .I (\syn181500/GROM ),
      .O (syn176960)
    );
    X_BUF \syn181500/XUSED (
      .I (\syn181500/FROM ),
      .O (syn181500)
    );
    defparam C18165.INIT = 16'hA05F;
    X_LUT4 C18165(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [23]),
      .ADR1 (VCC),
      .ADR2 (syn24500),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [23]),
      .O (\syn181501/GROM )
    );
    defparam C18164.INIT = 16'h9050;
    X_LUT4 C18164(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [24]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [24]),
      .ADR2 (syn176963),
      .ADR3 (syn24500),
      .O (\syn181501/FROM )
    );
    X_BUF \syn181501/YUSED (
      .I (\syn181501/GROM ),
      .O (syn176963)
    );
    X_BUF \syn181501/XUSED (
      .I (\syn181501/FROM ),
      .O (syn181501)
    );
    defparam C18163.INIT = 16'hA555;
    X_LUT4 C18163(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [21]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [21]),
      .ADR3 (syn24500),
      .O (\syn181502/GROM )
    );
    defparam C18162.INIT = 16'h9030;
    X_LUT4 C18162(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [22]),
      .ADR2 (syn176965),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [22]),
      .O (\syn181502/FROM )
    );
    X_BUF \syn181502/YUSED (
      .I (\syn181502/GROM ),
      .O (syn176965)
    );
    X_BUF \syn181502/XUSED (
      .I (\syn181502/FROM ),
      .O (syn181502)
    );
    defparam C18151.INIT = 16'h802A;
    X_LUT4 C18151(
      .ADR0 (syn176975),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [12]),
      .ADR2 (syn24500),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [12]),
      .O (\syn181522/GROM )
    );
    defparam C18150.INIT = 16'h8000;
    X_LUT4 C18150(
      .ADR0 (syn181506),
      .ADR1 (syn181504),
      .ADR2 (syn181507),
      .ADR3 (syn181505),
      .O (\syn181522/FROM )
    );
    X_BUF \syn181522/YUSED (
      .I (\syn181522/GROM ),
      .O (syn181507)
    );
    X_BUF \syn181522/XUSED (
      .I (\syn181522/FROM ),
      .O (syn181522)
    );
    defparam C18158.INIT = 16'hC03F;
    X_LUT4 C18158(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [17]),
      .ADR2 (syn24500),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [17]),
      .O (\syn181504/GROM )
    );
    defparam C18157.INIT = 16'h8070;
    X_LUT4 C18157(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [18]),
      .ADR2 (syn176969),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [18]),
      .O (\syn181504/FROM )
    );
    X_BUF \syn181504/YUSED (
      .I (\syn181504/GROM ),
      .O (syn176969)
    );
    X_BUF \syn181504/XUSED (
      .I (\syn181504/FROM ),
      .O (syn181504)
    );
    defparam C18156.INIT = 16'h9595;
    X_LUT4 C18156(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [15]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [15]),
      .ADR2 (syn24500),
      .ADR3 (VCC),
      .O (\syn181505/GROM )
    );
    defparam C18155.INIT = 16'h9030;
    X_LUT4 C18155(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [16]),
      .ADR2 (syn176971),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [16]),
      .O (\syn181505/FROM )
    );
    X_BUF \syn181505/YUSED (
      .I (\syn181505/GROM ),
      .O (syn176971)
    );
    X_BUF \syn181505/XUSED (
      .I (\syn181505/FROM ),
      .O (syn181505)
    );
    defparam C18154.INIT = 16'hA50F;
    X_LUT4 C18154(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [13]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_addr_out [13]),
      .ADR3 (syn24500),
      .O (\syn181506/GROM )
    );
    defparam C18153.INIT = 16'h9050;
    X_LUT4 C18153(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [14]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [14]),
      .ADR2 (syn176973),
      .ADR3 (syn24500),
      .O (\syn181506/FROM )
    );
    X_BUF \syn181506/YUSED (
      .I (\syn181506/GROM ),
      .O (syn176973)
    );
    X_BUF \syn181506/XUSED (
      .I (\syn181506/FROM ),
      .O (syn181506)
    );
    defparam C18149.INIT = 16'hA05F;
    X_LUT4 C18149(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [9]),
      .ADR1 (VCC),
      .ADR2 (syn24500),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [9]),
      .O (\syn181508/GROM )
    );
    defparam C18148.INIT = 16'h9030;
    X_LUT4 C18148(
      .ADR0 (syn24500),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [10]),
      .ADR2 (syn176977),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [10]),
      .O (\syn181508/FROM )
    );
    X_BUF \syn181508/YUSED (
      .I (\syn181508/GROM ),
      .O (syn176977)
    );
    X_BUF \syn181508/XUSED (
      .I (\syn181508/FROM ),
      .O (syn181508)
    );
    defparam C19351.INIT = 16'hCC00;
    X_LUT4 C19351(
      .ADR0 (VCC),
      .ADR1 (syn24500),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .O (\syn181510/GROM )
    );
    defparam C18146.INIT = 16'h2184;
    X_LUT4 C18146(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [5]),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_addr_out [6]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C104 ),
      .ADR3 (syn59978),
      .O (\syn181510/FROM )
    );
    X_BUF \syn181510/YUSED (
      .I (\syn181510/GROM ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C104 )
    );
    X_BUF \syn181510/XUSED (
      .I (\syn181510/FROM ),
      .O (syn181510)
    );
    defparam C17791.INIT = 16'hC000;
    X_LUT4 C17791(
      .ADR0 (VCC),
      .ADR1 (syn24519),
      .ADR2 (syn24524),
      .ADR3 (syn182355),
      .O (\N12544/GROM )
    );
    defparam C17790.INIT = 16'hFFF4;
    X_LUT4 C17790(
      .ADR0 (\bridge/pci_target_unit/del_sync/req_rty_exp_clr ),
      .ADR1 (\bridge/pci_target_unit/del_sync/req_rty_exp_reg ),
      .ADR2 (N12545),
      .ADR3 (\bridge/pci_target_unit/del_sync/req_comp_pending ),
      .O (\N12544/FROM )
    );
    X_BUF \N12544/YUSED (
      .I (\N12544/GROM ),
      .O (N12545)
    );
    X_BUF \N12544/XUSED (
      .I (\N12544/FROM ),
      .O (N12544)
    );
    defparam C19128.INIT = 16'hF8F0;
    X_LUT4 C19128(
      .ADR0 (syn24519),
      .ADR1 (syn17000),
      .ADR2 (syn19415),
      .ADR3 (syn24524),
      .O (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out/GROM )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_load_critical/C60 .INIT = 16'hF0FA;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_load_critical/C60 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/load_med_reg_w ),
      .ADR3 (N_IRDY),
      .O (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_sm_load_medium_reg_out/YUSED (
      .I (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out/GROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/load_med_reg_w )
    );
    X_BUF \bridge/pci_target_unit/pcit_sm_load_medium_reg_out/XUSED (
      .I (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out/FROM ),
      .O (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out )
    );
    defparam C19483.INIT = 16'h1111;
    X_LUT4 C19483(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [2]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [0]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn18863/GROM )
    );
    defparam C19478.INIT = 16'h3313;
    X_LUT4 C19478(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (syn17010),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .O (\syn18863/FROM )
    );
    X_BUF \syn18863/YUSED (
      .I (\syn18863/GROM ),
      .O (syn17010)
    );
    X_BUF \syn18863/XUSED (
      .I (\syn18863/FROM ),
      .O (syn18863)
    );
    defparam C19481.INIT = 16'h0FFF;
    X_LUT4 C19481(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .O (\syn18858/GROM )
    );
    defparam C19480.INIT = 16'h4090;
    X_LUT4 C19480(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [0]),
      .ADR1 (syn178535),
      .ADR2 (syn178547),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [2]),
      .O (\syn18858/FROM )
    );
    X_BUF \syn18858/YUSED (
      .I (\syn18858/GROM ),
      .O (syn178547)
    );
    X_BUF \syn18858/XUSED (
      .I (\syn18858/FROM ),
      .O (syn18858)
    );
    defparam C19984.INIT = 16'h2800;
    X_LUT4 C19984(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/del_completion_allow ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_bc_out [2]),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/map ),
      .ADR3 (\bridge/wishbone_slave_unit/wishbone_slave/del_addr_hit ),
      .O (\syn17669/GROM )
    );
    defparam C19983.INIT = 16'h9000;
    X_LUT4 C19983(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_bc_out [3]),
      .ADR1 (\bridge/wishbone_slave_unit/wbs_sm_del_bc_out [3]),
      .ADR2 (syn177332),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_bc_out [1]),
      .O (\syn17669/FROM )
    );
    X_BUF \syn17669/YUSED (
      .I (\syn17669/GROM ),
      .O (syn177332)
    );
    X_BUF \syn17669/XUSED (
      .I (\syn17669/FROM ),
      .O (syn17669)
    );
    defparam C19885.INIT = 16'h8888;
    X_LUT4 C19885(
      .ADR0 (\bridge/conf_pci_am1_out [18]),
      .ADR1 (\bridge/conf_pci_ba1_out [18]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn177570/GROM )
    );
    defparam C19884.INIT = 16'hEAC0;
    X_LUT4 C19884(
      .ADR0 (\bridge/configuration/C2318 ),
      .ADR1 (\bridge/configuration/C2360 ),
      .ADR2 (syn17051),
      .ADR3 (\bridge/configuration/wb_tran_addr1 [30]),
      .O (\syn177570/FROM )
    );
    X_BUF \syn177570/YUSED (
      .I (\syn177570/GROM ),
      .O (syn17051)
    );
    X_BUF \syn177570/XUSED (
      .I (\syn177570/FROM ),
      .O (syn177570)
    );
    defparam C19846.INIT = 16'hC0C0;
    X_LUT4 C19846(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_pci_ba1_out [16]),
      .ADR2 (\bridge/conf_pci_am1_out [16]),
      .ADR3 (VCC),
      .O (\syn177658/GROM )
    );
    defparam C19845.INIT = 16'hECA0;
    X_LUT4 C19845(
      .ADR0 (\bridge/configuration/C2360 ),
      .ADR1 (\bridge/configuration/wb_err_addr [28]),
      .ADR2 (syn17053),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn177658/FROM )
    );
    X_BUF \syn177658/YUSED (
      .I (\syn177658/GROM ),
      .O (syn17053)
    );
    X_BUF \syn177658/XUSED (
      .I (\syn177658/FROM ),
      .O (syn177658)
    );
    defparam C19796.INIT = 16'hF888;
    X_LUT4 C19796(
      .ADR0 (\bridge/conf_pci_ba0_out [13]),
      .ADR1 (\bridge/configuration/C2370 ),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [25]),
      .ADR3 (\bridge/configuration/C2318 ),
      .O (\syn177781/GROM )
    );
    defparam C19795.INIT = 16'hFFFE;
    X_LUT4 C19795(
      .ADR0 (syn177771),
      .ADR1 (syn18051),
      .ADR2 (syn177773),
      .ADR3 (syn177772),
      .O (\syn177781/FROM )
    );
    X_BUF \syn177781/YUSED (
      .I (\syn177781/GROM ),
      .O (syn177773)
    );
    X_BUF \syn177781/XUSED (
      .I (\syn177781/FROM ),
      .O (syn177781)
    );
    defparam C19740.INIT = 16'hF000;
    X_LUT4 C19740(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [21]),
      .ADR3 (\bridge/configuration/pci_base_addr1 [21]),
      .O (\syn177924/GROM )
    );
    defparam C19739.INIT = 16'hEAC0;
    X_LUT4 C19739(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/configuration/C2360 ),
      .ADR2 (syn17060),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [21]),
      .O (\syn177924/FROM )
    );
    X_BUF \syn177924/YUSED (
      .I (\syn177924/GROM ),
      .O (syn17060)
    );
    X_BUF \syn177924/XUSED (
      .I (\syn177924/FROM ),
      .O (syn177924)
    );
    defparam C19727.INIT = 16'hC0C0;
    X_LUT4 C19727(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_base_addr1 [20]),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [20]),
      .ADR3 (VCC),
      .O (\syn177957/GROM )
    );
    defparam C19726.INIT = 16'hEAC0;
    X_LUT4 C19726(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/configuration/C2360 ),
      .ADR2 (syn17061),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [20]),
      .O (\syn177957/FROM )
    );
    X_BUF \syn177957/YUSED (
      .I (\syn177957/GROM ),
      .O (syn17061)
    );
    X_BUF \syn177957/XUSED (
      .I (\syn177957/FROM ),
      .O (syn177957)
    );
    defparam C19688.INIT = 16'hCC00;
    X_LUT4 C19688(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_base_addr1 [17]),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [17]),
      .O (\syn178057/GROM )
    );
    defparam C19687.INIT = 16'hF888;
    X_LUT4 C19687(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [17]),
      .ADR2 (syn17064),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn178057/FROM )
    );
    X_BUF \syn178057/YUSED (
      .I (\syn178057/GROM ),
      .O (syn17064)
    );
    X_BUF \syn178057/XUSED (
      .I (\syn178057/FROM ),
      .O (syn178057)
    );
    defparam C19675.INIT = 16'hCC00;
    X_LUT4 C19675(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_base_addr1 [16]),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [16]),
      .O (\syn178095/GROM )
    );
    defparam C19674.INIT = 16'hF888;
    X_LUT4 C19674(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [16]),
      .ADR2 (syn17065),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn178095/FROM )
    );
    X_BUF \syn178095/YUSED (
      .I (\syn178095/GROM ),
      .O (syn17065)
    );
    X_BUF \syn178095/XUSED (
      .I (\syn178095/FROM ),
      .O (syn178095)
    );
    defparam C19616.INIT = 16'hAA00;
    X_LUT4 C19616(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [12]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/pci_base_addr1 [12]),
      .O (\syn178239/GROM )
    );
    defparam C19615.INIT = 16'hF888;
    X_LUT4 C19615(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [12]),
      .ADR2 (syn17070),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn178239/FROM )
    );
    X_BUF \syn178239/YUSED (
      .I (\syn178239/GROM ),
      .O (syn17070)
    );
    X_BUF \syn178239/XUSED (
      .I (\syn178239/FROM ),
      .O (syn178239)
    );
    defparam C19496.INIT = 16'hEAC0;
    X_LUT4 C19496(
      .ADR0 (\bridge/conf_pci_mem_io1_out ),
      .ADR1 (\bridge/configuration/C2304 ),
      .ADR2 (\bridge/configuration/wb_err_addr [0]),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn178522/GROM )
    );
    defparam C19495.INIT = 16'hFFFA;
    X_LUT4 C19495(
      .ADR0 (syn178514),
      .ADR1 (VCC),
      .ADR2 (syn178518),
      .ADR3 (syn178515),
      .O (\syn178522/FROM )
    );
    X_BUF \syn178522/YUSED (
      .I (\syn178522/GROM ),
      .O (syn178518)
    );
    X_BUF \syn178522/XUSED (
      .I (\syn178522/FROM ),
      .O (syn178522)
    );
    defparam C19394.INIT = 16'hECA0;
    X_LUT4 C19394(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .ADR1 (syn17086),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [4]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [4])
      ,
      .O (\bridge/wishbone_slave_unit/fifos/C3/N30/GROM )
    );
    defparam C19393.INIT = 16'hF8F8;
    X_LUT4 C19393(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [4]),
      .ADR1 (syn17087),
      .ADR2 (syn178727),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N30/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N30/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N30/GROM ),
      .O (syn178727)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N30/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N30/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N30 )
    );
    defparam C19401.INIT = 16'hFEFC;
    X_LUT4 C19401(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .ADR2 (syn60010),
      .ADR3 (syn19081),
      .O (\syn17087/GROM )
    );
    defparam C19399.INIT = 16'h3323;
    X_LUT4 C19399(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty ),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .ADR2 (syn19088),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty ),
      .O (\syn17087/FROM )
    );
    X_BUF \syn17087/YUSED (
      .I (\syn17087/GROM ),
      .O (syn19088)
    );
    X_BUF \syn17087/XUSED (
      .I (\syn17087/FROM ),
      .O (syn17087)
    );
    defparam C19406.INIT = 16'h0003;
    X_LUT4 C19406(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/err_recovery ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/cell8/GROM )
    );
    defparam C19405.INIT = 16'h0080;
    X_LUT4 C19405(
      .ADR0 (N12594),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_transaction_ready_out ),
      .ADR2 (syn178708),
      .ADR3 (\bridge/conf_wb_err_pending_out ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/cell8/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/cell8/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/cell8/GROM ),
      .O (syn178708)
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/cell8/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/cell8/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 )
    );
    defparam C19396.INIT = 16'hFFA0;
    X_LUT4 C19396(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/err_recovery ),
      .ADR1 (VCC),
      .ADR2 (N12594),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/cell8 ),
      .O (\syn17086/GROM )
    );
    defparam C19395.INIT = 16'h00A8;
    X_LUT4 C19395(
      .ADR0 (syn19075),
      .ADR1 (syn19085),
      .ADR2 (syn178718),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .O (\syn17086/FROM )
    );
    X_BUF \syn17086/YUSED (
      .I (\syn17086/GROM ),
      .O (syn178718)
    );
    X_BUF \syn17086/XUSED (
      .I (\syn17086/FROM ),
      .O (syn17086)
    );
    defparam C19392.INIT = 16'hECA0;
    X_LUT4 C19392(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [3])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .ADR2 (syn17086),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [3]),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N24/GROM )
    );
    defparam C19391.INIT = 16'hFCF0;
    X_LUT4 C19391(
      .ADR0 (VCC),
      .ADR1 (syn17087),
      .ADR2 (syn178732),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [3]),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N24/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N24/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N24/GROM ),
      .O (syn178732)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N24/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N24/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N24 )
    );
    defparam C19390.INIT = 16'hF888;
    X_LUT4 C19390(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [2]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [2])
      ,
      .ADR3 (syn17086),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N18/GROM )
    );
    defparam C19389.INIT = 16'hFAF0;
    X_LUT4 C19389(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [2]),
      .ADR1 (VCC),
      .ADR2 (syn178737),
      .ADR3 (syn17087),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N18/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N18/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N18/GROM ),
      .O (syn178737)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N18/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N18/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N18 )
    );
    defparam C19388.INIT = 16'hEAC0;
    X_LUT4 C19388(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [1])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [1]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .ADR3 (syn17086),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N12/GROM )
    );
    defparam C19387.INIT = 16'hFAF0;
    X_LUT4 C19387(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [1]),
      .ADR1 (VCC),
      .ADR2 (syn178742),
      .ADR3 (syn17087),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N12/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N12/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N12/GROM ),
      .O (syn178742)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N12/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N12/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N12 )
    );
    defparam C19386.INIT = 16'hEAC0;
    X_LUT4 C19386(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [0])
      ,
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [0]),
      .ADR3 (syn17086),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N6/GROM )
    );
    defparam C19385.INIT = 16'hF8F8;
    X_LUT4 C19385(
      .ADR0 (syn17087),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [0]),
      .ADR2 (syn178747),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N6/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N6/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N6/GROM ),
      .O (syn178747)
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N6/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N6/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N6 )
    );
    defparam C19314.INIT = 16'hFAAA;
    X_LUT4 C19314(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/state_backoff_reg ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .O (\syn19397/GROM )
    );
    defparam C19313.INIT = 16'hF200;
    X_LUT4 C19313(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/state_transfere_reg ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/disconect_wo_data_reg ),
      .ADR2 (syn178873),
      .ADR3 (syn16919),
      .O (\syn19397/FROM )
    );
    X_BUF \syn19397/YUSED (
      .I (\syn19397/GROM ),
      .O (syn178873)
    );
    X_BUF \syn19397/XUSED (
      .I (\syn19397/FROM ),
      .O (syn19397)
    );
    defparam C19248.INIT = 16'hAA0C;
    X_LUT4 C19248(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_raddr [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .O (\bridge/pci_target_unit/fifos/C10/N30/GROM )
    );
    defparam C19247.INIT = 16'hF0F8;
    X_LUT4 C19247(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_raddr_0 [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR2 (syn179034),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .O (\bridge/pci_target_unit/fifos/C10/N30/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N30/YUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N30/GROM ),
      .O (syn179034)
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N30/XUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N30/FROM ),
      .O (\bridge/pci_target_unit/fifos/C10/N30 )
    );
    defparam C19262.INIT = 16'hC0C0;
    X_LUT4 C19262(
      .ADR0 (VCC),
      .ADR1 (syn178999),
      .ADR2 (syn178998),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[1]/GROM )
    );
    defparam C19261.INIT = 16'h80A8;
    X_LUT4 C19261(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .ADR1 (ERR_I),
      .ADR2 (syn19555),
      .ADR3 (ACK_I),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[1]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out<1>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[1]/GROM ),
      .O (syn19555)
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out<1>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[1]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out [1])
    );
    defparam C19245.INIT = 16'hBA10;
    X_LUT4 C19245(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_raddr [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_waddr [3]),
      .O (\bridge/pci_target_unit/fifos/C10/N24/GROM )
    );
    defparam C19244.INIT = 16'hF4F0;
    X_LUT4 C19244(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR2 (syn179042),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_raddr_0 [3]),
      .O (\bridge/pci_target_unit/fifos/C10/N24/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N24/YUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N24/GROM ),
      .O (syn179042)
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N24/XUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N24/FROM ),
      .O (\bridge/pci_target_unit/fifos/C10/N24 )
    );
    defparam C19242.INIT = 16'hDC10;
    X_LUT4 C19242(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_raddr [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_waddr [2]),
      .O (\bridge/pci_target_unit/fifos/C10/N18/GROM )
    );
    defparam C19241.INIT = 16'hF2F0;
    X_LUT4 C19241(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .ADR2 (syn179050),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_raddr_0 [2]),
      .O (\bridge/pci_target_unit/fifos/C10/N18/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N18/YUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N18/GROM ),
      .O (syn179050)
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N18/XUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N18/FROM ),
      .O (\bridge/pci_target_unit/fifos/C10/N18 )
    );
    defparam C19239.INIT = 16'h8B88;
    X_LUT4 C19239(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [1]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_raddr [1]),
      .O (\bridge/pci_target_unit/fifos/C10/N12/GROM )
    );
    defparam C19238.INIT = 16'hF4F0;
    X_LUT4 C19238(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_raddr_0 [1]),
      .ADR2 (syn179058),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .O (\bridge/pci_target_unit/fifos/C10/N12/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N12/YUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N12/GROM ),
      .O (syn179058)
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N12/XUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N12/FROM ),
      .O (\bridge/pci_target_unit/fifos/C10/N12 )
    );
    defparam C19236.INIT = 16'hAA0C;
    X_LUT4 C19236(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_raddr [0]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .O (\bridge/pci_target_unit/fifos/C10/N6/GROM )
    );
    defparam C19235.INIT = 16'hF2F0;
    X_LUT4 C19235(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .ADR2 (syn179066),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_raddr_0 [0]),
      .O (\bridge/pci_target_unit/fifos/C10/N6/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N6/YUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N6/GROM ),
      .O (syn179066)
    );
    X_BUF \bridge/pci_target_unit/fifos/C10/N6/XUSED (
      .I (\bridge/pci_target_unit/fifos/C10/N6/FROM ),
      .O (\bridge/pci_target_unit/fifos/C10/N6 )
    );
    defparam C19217.INIT = 16'h0404;
    X_LUT4 C19217(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_full ),
      .ADR2 (\bridge/pci_target_unit/fifos_pciw_full_out ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/in_count_en/GROM )
    );
    defparam C17935.INIT = 16'h3230;
    X_LUT4 C17935(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR1 (N12616),
      .ADR2 (syn19671),
      .ADR3 (\bridge/in_reg_frame_out ),
      .O (\bridge/pci_target_unit/fifos/in_count_en/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/in_count_en/YUSED (
      .I (\bridge/pci_target_unit/fifos/in_count_en/GROM ),
      .O (syn19671)
    );
    X_BUF \bridge/pci_target_unit/fifos/in_count_en/XUSED (
      .I (\bridge/pci_target_unit/fifos/in_count_en/FROM ),
      .O (\bridge/pci_target_unit/fifos/in_count_en )
    );
    defparam C19141.INIT = 16'hFF05;
    X_LUT4 C19141(
      .ADR0 (\bridge/pci_target_unit/pcit_if_pcir_fifo_data_err_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR3 (\bridge/in_reg_irdy_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm/GROM )
    );
    defparam C19140.INIT = 16'hC4C4;
    X_LUT4 C19140(
      .ADR0 (\bridge/pci_target_unit/pcit_if_disconect_wo_data_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/N64 ),
      .ADR2 (syn179294),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/trdy_w_frm/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm/GROM ),
      .O (syn179294)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/trdy_w_frm/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm )
    );
    defparam C18867.INIT = 16'h80A0;
    X_LUT4 C18867(
      .ADR0 (syn20406),
      .ADR1 (syn20373),
      .ADR2 (syn179711),
      .ADR3 (\bridge/pciu_conf_offset_out [2]),
      .O (\bridge/configuration/C285/N34/GROM )
    );
    defparam C18866.INIT = 16'h00F0;
    X_LUT4 C18866(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn17097),
      .ADR3 (\bridge/in_reg_cbe_out [3]),
      .O (\bridge/configuration/C285/N34/FROM )
    );
    X_BUF \bridge/configuration/C285/N34/YUSED (
      .I (\bridge/configuration/C285/N34/GROM ),
      .O (syn17097)
    );
    X_BUF \bridge/configuration/C285/N34/XUSED (
      .I (\bridge/configuration/C285/N34/FROM ),
      .O (\bridge/configuration/C285/N34 )
    );
    defparam C18885.INIT = 16'hF8F0;
    X_LUT4 C18885(
      .ADR0 (syn179694),
      .ADR1 (syn20371),
      .ADR2 (\bridge/pciu_conf_offset_out [2]),
      .ADR3 (syn20360),
      .O (\syn20406/GROM )
    );
    defparam C18883.INIT = 16'h64A0;
    X_LUT4 C18883(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (syn60090),
      .ADR2 (syn20389),
      .ADR3 (syn60111),
      .O (\syn20406/FROM )
    );
    X_BUF \syn20406/YUSED (
      .I (\syn20406/GROM ),
      .O (syn20389)
    );
    X_BUF \syn20406/XUSED (
      .I (\syn20406/FROM ),
      .O (syn20406)
    );
    defparam C18912.INIT = 16'h000F;
    X_LUT4 C18912(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pciu_conf_offset_out [7]),
      .ADR3 (\bridge/pciu_conf_offset_out [6]),
      .O (\syn20371/GROM )
    );
    defparam C18892.INIT = 16'h31FF;
    X_LUT4 C18892(
      .ADR0 (\bridge/pciu_conf_offset_out [3]),
      .ADR1 (\bridge/pciu_conf_offset_out [5]),
      .ADR2 (syn60111),
      .ADR3 (\bridge/pciu_conf_offset_out [4]),
      .O (\syn20371/FROM )
    );
    X_BUF \syn20371/YUSED (
      .I (\syn20371/GROM ),
      .O (syn60111)
    );
    X_BUF \syn20371/XUSED (
      .I (\syn20371/FROM ),
      .O (syn20371)
    );
    defparam C18887.INIT = 16'hDDFC;
    X_LUT4 C18887(
      .ADR0 (\bridge/pciu_conf_offset_out [3]),
      .ADR1 (\bridge/pciu_conf_offset_out [4]),
      .ADR2 (\bridge/pciu_conf_offset_out [7]),
      .ADR3 (\bridge/pciu_conf_offset_out [6]),
      .O (\syn179694/GROM )
    );
    defparam C18886.INIT = 16'hF030;
    X_LUT4 C18886(
      .ADR0 (VCC),
      .ADR1 (\bridge/pciu_conf_offset_out [5]),
      .ADR2 (syn20359),
      .ADR3 (\bridge/pciu_conf_offset_out [6]),
      .O (\syn179694/FROM )
    );
    X_BUF \syn179694/YUSED (
      .I (\syn179694/GROM ),
      .O (syn20359)
    );
    X_BUF \syn179694/XUSED (
      .I (\syn179694/FROM ),
      .O (syn179694)
    );
    defparam C18873.INIT = 16'h0001;
    X_LUT4 C18873(
      .ADR0 (\bridge/configuration/C1973 ),
      .ADR1 (\bridge/configuration/C1959 ),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/configuration/C1955 ),
      .O (\syn179711/GROM )
    );
    defparam C18868.INIT = 16'h8080;
    X_LUT4 C18868(
      .ADR0 (syn179707),
      .ADR1 (syn179709),
      .ADR2 (syn179708),
      .ADR3 (VCC),
      .O (\syn179711/FROM )
    );
    X_BUF \syn179711/YUSED (
      .I (\syn179711/GROM ),
      .O (syn179708)
    );
    X_BUF \syn179711/XUSED (
      .I (\syn179711/FROM ),
      .O (syn179711)
    );
    defparam C18880.INIT = 16'h2020;
    X_LUT4 C18880(
      .ADR0 (\bridge/pciu_conf_offset_out [7]),
      .ADR1 (\bridge/pciu_conf_offset_out [6]),
      .ADR2 (syn60090),
      .ADR3 (VCC),
      .O (\syn179707/GROM )
    );
    defparam C18879.INIT = 16'h0001;
    X_LUT4 C18879(
      .ADR0 (\bridge/configuration/C1941 ),
      .ADR1 (\bridge/configuration/C1925 ),
      .ADR2 (\bridge/configuration/C1951 ),
      .ADR3 (\bridge/configuration/C1929 ),
      .O (\syn179707/FROM )
    );
    X_BUF \syn179707/YUSED (
      .I (\syn179707/GROM ),
      .O (\bridge/configuration/C1951 )
    );
    X_BUF \syn179707/XUSED (
      .I (\syn179707/FROM ),
      .O (syn179707)
    );
    defparam C18911.INIT = 16'h0055;
    X_LUT4 C18911(
      .ADR0 (\bridge/pciu_conf_offset_out [4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pciu_conf_offset_out [5]),
      .O (\bridge/configuration/C1959/GROM )
    );
    defparam C18876.INIT = 16'h2000;
    X_LUT4 C18876(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (syn179659),
      .ADR3 (syn17004),
      .O (\bridge/configuration/C1959/FROM )
    );
    X_BUF \bridge/configuration/C1959/YUSED (
      .I (\bridge/configuration/C1959/GROM ),
      .O (syn179659)
    );
    X_BUF \bridge/configuration/C1959/XUSED (
      .I (\bridge/configuration/C1959/FROM ),
      .O (\bridge/configuration/C1959 )
    );
    defparam C18917.INIT = 16'h2000;
    X_LUT4 C18917(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR1 (syn19366),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/state_transfere_reg ),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .O (\syn179709/GROM )
    );
    defparam C18869.INIT = 16'h0010;
    X_LUT4 C18869(
      .ADR0 (\bridge/configuration/C1987 ),
      .ADR1 (syn60110),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/configuration/C1989 ),
      .O (\syn179709/FROM )
    );
    X_BUF \syn179709/YUSED (
      .I (\syn179709/GROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 )
    );
    X_BUF \syn179709/XUSED (
      .I (\syn179709/FROM ),
      .O (syn179709)
    );
    defparam C18787.INIT = 16'hCC00;
    X_LUT4 C18787(
      .ADR0 (VCC),
      .ADR1 (syn16916),
      .ADR2 (VCC),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn20486/GROM )
    );
    defparam C18786.INIT = 16'hF0E0;
    X_LUT4 C18786(
      .ADR0 (syn179850),
      .ADR1 (syn179855),
      .ADR2 (syn181260),
      .ADR3 (syn179851),
      .O (\syn20486/FROM )
    );
    X_BUF \syn20486/YUSED (
      .I (\syn20486/GROM ),
      .O (syn181260)
    );
    X_BUF \syn20486/XUSED (
      .I (\syn20486/FROM ),
      .O (syn20486)
    );
    defparam C18790.INIT = 16'hEAC0;
    X_LUT4 C18790(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/configuration/wb_img_ctrl1[0] ),
      .ADR2 (\bridge/configuration/C1959 ),
      .ADR3 (\bridge/conf_wb_mem_io1_out ),
      .O (\syn179855/GROM )
    );
    defparam C18789.INIT = 16'hFFFE;
    X_LUT4 C18789(
      .ADR0 (syn179846),
      .ADR1 (syn179848),
      .ADR2 (syn179849),
      .ADR3 (syn179847),
      .O (\syn179855/FROM )
    );
    X_BUF \syn179855/YUSED (
      .I (\syn179855/GROM ),
      .O (syn179849)
    );
    X_BUF \syn179855/XUSED (
      .I (\syn179855/FROM ),
      .O (syn179855)
    );
    defparam C18881.INIT = 16'h8000;
    X_LUT4 C18881(
      .ADR0 (syn17002),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (\bridge/pciu_conf_offset_out [7]),
      .ADR3 (\bridge/pciu_conf_offset_out [2]),
      .O (\syn179846/GROM )
    );
    defparam C18795.INIT = 16'hC0C0;
    X_LUT4 C18795(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/int_prop_en ),
      .ADR2 (\bridge/configuration/C1925 ),
      .ADR3 (VCC),
      .O (\syn179846/FROM )
    );
    X_BUF \syn179846/YUSED (
      .I (\syn179846/GROM ),
      .O (\bridge/configuration/C1925 )
    );
    X_BUF \syn179846/XUSED (
      .I (\syn179846/FROM ),
      .O (syn179846)
    );
    defparam C18782.INIT = 16'hECA0;
    X_LUT4 C18782(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [0]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_data_out [0]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (syn20493),
      .O (\syn20502/GROM )
    );
    defparam C18781.INIT = 16'h5450;
    X_LUT4 C18781(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn179869),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [0]),
      .O (\syn20502/FROM )
    );
    X_BUF \syn20502/YUSED (
      .I (\syn20502/GROM ),
      .O (syn179869)
    );
    X_BUF \syn20502/XUSED (
      .I (\syn20502/FROM ),
      .O (syn20502)
    );
    defparam C18784.INIT = 16'h8080;
    X_LUT4 C18784(
      .ADR0 (syn18858),
      .ADR1 (syn20490),
      .ADR2 (syn18863),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C155/GROM )
    );
    defparam C18783.INIT = 16'h0505;
    X_LUT4 C18783(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (VCC),
      .ADR2 (syn20493),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C155/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/C155/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C155/GROM ),
      .O (syn20493)
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/C155/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C155/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 )
    );
    defparam C18776.INIT = 16'h8800;
    X_LUT4 C18776(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/conf_io_space_enable_out ),
      .ADR2 (VCC),
      .ADR3 (syn17098),
      .O (\syn179882/GROM )
    );
    defparam C18773.INIT = 16'hFEFA;
    X_LUT4 C18773(
      .ADR0 (syn20484),
      .ADR1 (syn17120),
      .ADR2 (syn20482),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn179882/FROM )
    );
    X_BUF \syn179882/YUSED (
      .I (\syn179882/GROM ),
      .O (syn20482)
    );
    X_BUF \syn179882/XUSED (
      .I (\syn179882/FROM ),
      .O (syn179882)
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_sm/ad_iob_ce/C34 .INIT = 16'hAEAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_sm/ad_iob_ce/C34 (
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/load_force ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (N_TRDY),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_bc_out [0]),
      .O (\bridge/output_backup/data_load/GROM )
    );
    defparam C18760.INIT = 16'hFFF0;
    X_LUT4 C18760(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_mux_mas_load_in ),
      .ADR3 (\bridge/pci_mux_tar_load_in ),
      .O (\bridge/output_backup/data_load/FROM )
    );
    X_BUF \bridge/output_backup/data_load/YUSED (
      .I (\bridge/output_backup/data_load/GROM ),
      .O (\bridge/pci_mux_mas_load_in )
    );
    X_BUF \bridge/output_backup/data_load/XUSED (
      .I (\bridge/output_backup/data_load/FROM ),
      .O (\bridge/output_backup/data_load )
    );
    defparam C18751.INIT = 16'hF888;
    X_LUT4 C18751(
      .ADR0 (syn17104),
      .ADR1 (\bridge/configuration/interrupt_line [1]),
      .ADR2 (syn17101),
      .ADR3 (\bridge/conf_cache_line_size_out [1]),
      .O (\syn20532/GROM )
    );
    defparam C18750.INIT = 16'hFEFC;
    X_LUT4 C18750(
      .ADR0 (syn20523),
      .ADR1 (syn179919),
      .ADR2 (syn179920),
      .ADR3 (syn16916),
      .O (\syn20532/FROM )
    );
    X_BUF \syn20532/YUSED (
      .I (\syn20532/GROM ),
      .O (syn179920)
    );
    X_BUF \syn20532/XUSED (
      .I (\syn20532/FROM ),
      .O (syn20532)
    );
    defparam C18755.INIT = 16'hECA0;
    X_LUT4 C18755(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/configuration/C1967 ),
      .ADR2 (\bridge/configuration/pci_err_addr [1]),
      .ADR3 (\bridge/configuration/pci_err_data [1]),
      .O (\syn20523/GROM )
    );
    defparam C18754.INIT = 16'hFFFE;
    X_LUT4 C18754(
      .ADR0 (syn179912),
      .ADR1 (syn179910),
      .ADR2 (syn179913),
      .ADR3 (syn179911),
      .O (\syn20523/FROM )
    );
    X_BUF \syn20523/YUSED (
      .I (\syn20523/GROM ),
      .O (syn179913)
    );
    X_BUF \syn20523/XUSED (
      .I (\syn20523/FROM ),
      .O (syn20523)
    );
    defparam C18753.INIT = 16'hA280;
    X_LUT4 C18753(
      .ADR0 (syn19366),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [1]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [1]),
      .O (\syn179919/GROM )
    );
    defparam C18752.INIT = 16'hFAF0;
    X_LUT4 C18752(
      .ADR0 (syn17098),
      .ADR1 (VCC),
      .ADR2 (syn179918),
      .ADR3 (\bridge/conf_mem_space_enable_out ),
      .O (\syn179919/FROM )
    );
    X_BUF \syn179919/YUSED (
      .I (\syn179919/GROM ),
      .O (syn179918)
    );
    X_BUF \syn179919/XUSED (
      .I (\syn179919/FROM ),
      .O (syn179919)
    );
    defparam C18741.INIT = 16'hFEFC;
    X_LUT4 C18741(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (syn179948),
      .ADR2 (syn179951),
      .ADR3 (\bridge/configuration/pci_err_addr [2]),
      .O (\syn20564/GROM )
    );
    defparam C18740.INIT = 16'hFE00;
    X_LUT4 C18740(
      .ADR0 (syn179950),
      .ADR1 (syn179949),
      .ADR2 (syn179954),
      .ADR3 (syn16916),
      .O (\syn20564/FROM )
    );
    X_BUF \syn20564/YUSED (
      .I (\syn20564/GROM ),
      .O (syn179954)
    );
    X_BUF \syn20564/XUSED (
      .I (\syn20564/FROM ),
      .O (syn20564)
    );
    defparam C18736.INIT = 16'hF888;
    X_LUT4 C18736(
      .ADR0 (\bridge/configuration/interrupt_line [2]),
      .ADR1 (syn17104),
      .ADR2 (syn17101),
      .ADR3 (\bridge/conf_cache_line_size_out [2]),
      .O (\syn179960/GROM )
    );
    defparam C18735.INIT = 16'hFEFC;
    X_LUT4 C18735(
      .ADR0 (\bridge/conf_pci_master_enable_out ),
      .ADR1 (syn179957),
      .ADR2 (syn179959),
      .ADR3 (syn17098),
      .O (\syn179960/FROM )
    );
    X_BUF \syn179960/YUSED (
      .I (\syn179960/GROM ),
      .O (syn179959)
    );
    X_BUF \syn179960/XUSED (
      .I (\syn179960/FROM ),
      .O (syn179960)
    );
    defparam C18721.INIT = 16'hFF80;
    X_LUT4 C18721(
      .ADR0 (\bridge/configuration/pci_err_addr [3]),
      .ADR1 (\bridge/configuration/C1971 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (syn179985),
      .O (\syn20598/GROM )
    );
    defparam C18720.INIT = 16'hFFFE;
    X_LUT4 C18720(
      .ADR0 (syn179988),
      .ADR1 (syn179987),
      .ADR2 (syn179989),
      .ADR3 (syn179986),
      .O (\syn20598/FROM )
    );
    X_BUF \syn20598/YUSED (
      .I (\syn20598/GROM ),
      .O (syn179989)
    );
    X_BUF \syn20598/XUSED (
      .I (\syn20598/FROM ),
      .O (syn20598)
    );
    defparam C18719.INIT = 16'hF888;
    X_LUT4 C18719(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_data_out [3]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [3]),
      .O (\syn20611/GROM )
    );
    defparam C18718.INIT = 16'h3230;
    X_LUT4 C18718(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180000),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [3]),
      .O (\syn20611/FROM )
    );
    X_BUF \syn20611/YUSED (
      .I (\syn20611/GROM ),
      .O (syn180000)
    );
    X_BUF \syn20611/XUSED (
      .I (\syn20611/FROM ),
      .O (syn20611)
    );
    defparam C18705.INIT = 16'hECA0;
    X_LUT4 C18705(
      .ADR0 (\bridge/conf_cache_line_size_out [4]),
      .ADR1 (syn17104),
      .ADR2 (syn17101),
      .ADR3 (\bridge/configuration/interrupt_line [4]),
      .O (\syn20635/GROM )
    );
    defparam C18704.INIT = 16'hFFFE;
    X_LUT4 C18704(
      .ADR0 (syn180031),
      .ADR1 (syn180032),
      .ADR2 (syn180033),
      .ADR3 (syn180030),
      .O (\syn20635/FROM )
    );
    X_BUF \syn20635/YUSED (
      .I (\syn20635/GROM ),
      .O (syn180033)
    );
    X_BUF \syn20635/XUSED (
      .I (\syn20635/FROM ),
      .O (syn20635)
    );
    defparam C18710.INIT = 16'hCC00;
    X_LUT4 C18710(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/C1935 ),
      .ADR2 (VCC),
      .ADR3 (syn16916),
      .O (\syn180031/GROM )
    );
    defparam C18709.INIT = 16'hEAC0;
    X_LUT4 C18709(
      .ADR0 (\bridge/configuration/wb_err_addr [4]),
      .ADR1 (\bridge/configuration/wb_err_data [4]),
      .ADR2 (syn17111),
      .ADR3 (syn17110),
      .O (\syn180031/FROM )
    );
    X_BUF \syn180031/YUSED (
      .I (\syn180031/GROM ),
      .O (syn17111)
    );
    X_BUF \syn180031/XUSED (
      .I (\syn180031/FROM ),
      .O (syn180031)
    );
    defparam C18788.INIT = 16'h0010;
    X_LUT4 C18788(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR1 (syn19366),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/out_bckp_devsel_out ),
      .O (\syn17110/GROM )
    );
    defparam C18711.INIT = 16'hC0C0;
    X_LUT4 C18711(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/C1937 ),
      .ADR2 (syn16916),
      .ADR3 (VCC),
      .O (\syn17110/FROM )
    );
    X_BUF \syn17110/YUSED (
      .I (\syn17110/GROM ),
      .O (syn16916)
    );
    X_BUF \syn17110/XUSED (
      .I (\syn17110/FROM ),
      .O (syn17110)
    );
    defparam C18707.INIT = 16'hC0C0;
    X_LUT4 C18707(
      .ADR0 (VCC),
      .ADR1 (syn16916),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (VCC),
      .O (\syn180032/GROM )
    );
    defparam C18706.INIT = 16'hEAC0;
    X_LUT4 C18706(
      .ADR0 (syn17107),
      .ADR1 (\bridge/configuration/pci_err_data [4]),
      .ADR2 (syn17109),
      .ADR3 (\bridge/configuration/pci_err_addr [4]),
      .O (\syn180032/FROM )
    );
    X_BUF \syn180032/YUSED (
      .I (\syn180032/GROM ),
      .O (syn17109)
    );
    X_BUF \syn180032/XUSED (
      .I (\syn180032/FROM ),
      .O (syn180032)
    );
    defparam C18692.INIT = 16'hECA0;
    X_LUT4 C18692(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_data_out [5]),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [5]),
      .O (\syn20672/GROM )
    );
    defparam C18691.INIT = 16'h3230;
    X_LUT4 C18691(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [5]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180064),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\syn20672/FROM )
    );
    X_BUF \syn20672/YUSED (
      .I (\syn20672/GROM ),
      .O (syn180064)
    );
    X_BUF \syn20672/XUSED (
      .I (\syn20672/FROM ),
      .O (syn20672)
    );
    defparam C18684.INIT = 16'hEAC0;
    X_LUT4 C18684(
      .ADR0 (\bridge/configuration/pci_err_data [6]),
      .ADR1 (syn16983),
      .ADR2 (\bridge/configuration/pci_err_addr [6]),
      .ADR3 (syn16985),
      .O (\syn20688/GROM )
    );
    defparam C18683.INIT = 16'hFFFE;
    X_LUT4 C18683(
      .ADR0 (syn180082),
      .ADR1 (syn180083),
      .ADR2 (syn180084),
      .ADR3 (syn180081),
      .O (\syn20688/FROM )
    );
    X_BUF \syn20688/YUSED (
      .I (\syn20688/GROM ),
      .O (syn180084)
    );
    X_BUF \syn20688/XUSED (
      .I (\syn20688/FROM ),
      .O (syn20688)
    );
    defparam C18909.INIT = 16'h4444;
    X_LUT4 C18909(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/configuration/C2003 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn180082/GROM )
    );
    defparam C18686.INIT = 16'hF888;
    X_LUT4 C18686(
      .ADR0 (\bridge/configuration/config_addr[6] ),
      .ADR1 (syn17016),
      .ADR2 (syn17099),
      .ADR3 (\bridge/conf_perr_response_out ),
      .O (\syn180082/FROM )
    );
    X_BUF \syn180082/YUSED (
      .I (\syn180082/GROM ),
      .O (syn17099)
    );
    X_BUF \syn180082/XUSED (
      .I (\syn180082/FROM ),
      .O (syn180082)
    );
    defparam C18682.INIT = 16'hF888;
    X_LUT4 C18682(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [6]),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [6]),
      .O (\syn20701/GROM )
    );
    defparam C18681.INIT = 16'h3230;
    X_LUT4 C18681(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [6]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180095),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\syn20701/FROM )
    );
    X_BUF \syn20701/YUSED (
      .I (\syn20701/GROM ),
      .O (syn180095)
    );
    X_BUF \syn20701/XUSED (
      .I (\syn20701/FROM ),
      .O (syn20701)
    );
    defparam C18673.INIT = 16'hECA0;
    X_LUT4 C18673(
      .ADR0 (\bridge/configuration/interrupt_line [7]),
      .ADR1 (\bridge/conf_cache_line_size_out [7]),
      .ADR2 (syn17104),
      .ADR3 (syn17101),
      .O (\syn20720/GROM )
    );
    defparam C18672.INIT = 16'hFFFE;
    X_LUT4 C18672(
      .ADR0 (syn180121),
      .ADR1 (syn180122),
      .ADR2 (syn180123),
      .ADR3 (syn180120),
      .O (\syn20720/FROM )
    );
    X_BUF \syn20720/YUSED (
      .I (\syn20720/GROM ),
      .O (syn180123)
    );
    X_BUF \syn20720/XUSED (
      .I (\syn20720/FROM ),
      .O (syn20720)
    );
    defparam C18667.INIT = 16'hF888;
    X_LUT4 C18667(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [8]),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [8]),
      .O (\syn20759/GROM )
    );
    defparam C18666.INIT = 16'h5450;
    X_LUT4 C18666(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn180167),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [8]),
      .O (\syn20759/FROM )
    );
    X_BUF \syn20759/YUSED (
      .I (\syn20759/GROM ),
      .O (syn180167)
    );
    X_BUF \syn20759/XUSED (
      .I (\syn20759/FROM ),
      .O (syn20759)
    );
    defparam C18657.INIT = 16'h8800;
    X_LUT4 C18657(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn17102),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_latency_tim_out [0]),
      .O (\syn180176/GROM )
    );
    defparam C18656.INIT = 16'hC8C8;
    X_LUT4 C18656(
      .ADR0 (syn180138),
      .ADR1 (syn60038),
      .ADR2 (syn180141),
      .ADR3 (VCC),
      .O (\syn180176/FROM )
    );
    X_BUF \syn180176/YUSED (
      .I (\syn180176/GROM ),
      .O (syn180141)
    );
    X_BUF \syn180176/XUSED (
      .I (\syn180176/FROM ),
      .O (syn180176)
    );
    defparam C18640.INIT = 16'hFFFE;
    X_LUT4 C18640(
      .ADR0 (syn20773),
      .ADR1 (syn20772),
      .ADR2 (syn20771),
      .ADR3 (syn20770),
      .O (\syn137911/GROM )
    );
    defparam C18639.INIT = 16'hFFFE;
    X_LUT4 C18639(
      .ADR0 (syn17121),
      .ADR1 (syn180205),
      .ADR2 (syn180209),
      .ADR3 (syn17017),
      .O (\syn137911/FROM )
    );
    X_BUF \syn137911/YUSED (
      .I (\syn137911/GROM ),
      .O (syn180209)
    );
    X_BUF \syn137911/XUSED (
      .I (\syn137911/FROM ),
      .O (syn137911)
    );
    defparam C18636.INIT = 16'hFFFE;
    X_LUT4 C18636(
      .ADR0 (syn20770),
      .ADR1 (syn20769),
      .ADR2 (syn20772),
      .ADR3 (syn20771),
      .O (\syn180212/GROM )
    );
    defparam C18635.INIT = 16'hAAA8;
    X_LUT4 C18635(
      .ADR0 (syn180250),
      .ADR1 (syn20773),
      .ADR2 (syn180202),
      .ADR3 (syn180198),
      .O (\syn180212/FROM )
    );
    X_BUF \syn180212/YUSED (
      .I (\syn180212/GROM ),
      .O (syn180202)
    );
    X_BUF \syn180212/XUSED (
      .I (\syn180212/FROM ),
      .O (syn180212)
    );
    defparam C18623.INIT = 16'hF888;
    X_LUT4 C18623(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [10]),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [10]),
      .O (\syn20817/GROM )
    );
    defparam C18622.INIT = 16'h00F8;
    X_LUT4 C18622(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [10]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn180258),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn20817/FROM )
    );
    X_BUF \syn20817/YUSED (
      .I (\syn20817/GROM ),
      .O (syn180258)
    );
    X_BUF \syn20817/XUSED (
      .I (\syn20817/FROM ),
      .O (syn20817)
    );
    defparam C18614.INIT = 16'hFCCC;
    X_LUT4 C18614(
      .ADR0 (VCC),
      .ADR1 (syn180282),
      .ADR2 (syn17101),
      .ADR3 (\bridge/conf_latency_tim_out [3]),
      .O (\syn20835/GROM )
    );
    defparam C18613.INIT = 16'hFFFC;
    X_LUT4 C18613(
      .ADR0 (VCC),
      .ADR1 (syn180284),
      .ADR2 (syn180285),
      .ADR3 (syn180283),
      .O (\syn20835/FROM )
    );
    X_BUF \syn20835/YUSED (
      .I (\syn20835/GROM ),
      .O (syn180285)
    );
    X_BUF \syn20835/XUSED (
      .I (\syn20835/FROM ),
      .O (syn20835)
    );
    defparam C18616.INIT = 16'hA280;
    X_LUT4 C18616(
      .ADR0 (syn19366),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [11]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [11]),
      .O (\syn180282/GROM )
    );
    defparam C18615.INIT = 16'hF8F0;
    X_LUT4 C18615(
      .ADR0 (\bridge/configuration/C1929 ),
      .ADR1 (\bridge/configuration/config_addr[11] ),
      .ADR2 (syn180281),
      .ADR3 (syn16916),
      .O (\syn180282/FROM )
    );
    X_BUF \syn180282/YUSED (
      .I (\syn180282/GROM ),
      .O (syn180281)
    );
    X_BUF \syn180282/XUSED (
      .I (\syn180282/FROM ),
      .O (syn180282)
    );
    defparam C18607.INIT = 16'hECCC;
    X_LUT4 C18607(
      .ADR0 (syn60110),
      .ADR1 (\bridge/configuration/C2001 ),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [12]),
      .ADR3 (\bridge/configuration/pci_base_addr1 [12]),
      .O (\syn180321/GROM )
    );
    defparam C18606.INIT = 16'hFFF8;
    X_LUT4 C18606(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/configuration/pci_err_addr [12]),
      .ADR2 (syn180313),
      .ADR3 (syn20853),
      .O (\syn180321/FROM )
    );
    X_BUF \syn180321/YUSED (
      .I (\syn180321/GROM ),
      .O (syn180313)
    );
    X_BUF \syn180321/XUSED (
      .I (\syn180321/FROM ),
      .O (syn180321)
    );
    defparam C18602.INIT = 16'hEAC0;
    X_LUT4 C18602(
      .ADR0 (\bridge/configuration/pci_err_data [12]),
      .ADR1 (\bridge/configuration/C1937 ),
      .ADR2 (\bridge/configuration/wb_err_addr [12]),
      .ADR3 (\bridge/configuration/C1967 ),
      .O (\syn180322/GROM )
    );
    defparam C18601.INIT = 16'hFFFE;
    X_LUT4 C18601(
      .ADR0 (syn180315),
      .ADR1 (syn180316),
      .ADR2 (syn180317),
      .ADR3 (syn180314),
      .O (\syn180322/FROM )
    );
    X_BUF \syn180322/YUSED (
      .I (\syn180322/GROM ),
      .O (syn180317)
    );
    X_BUF \syn180322/XUSED (
      .I (\syn180322/FROM ),
      .O (syn180322)
    );
    defparam C18599.INIT = 16'hECA0;
    X_LUT4 C18599(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [12]),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [12]),
      .O (\syn20882/GROM )
    );
    defparam C18598.INIT = 16'h3230;
    X_LUT4 C18598(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [12]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180329),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\syn20882/FROM )
    );
    X_BUF \syn20882/YUSED (
      .I (\syn20882/GROM ),
      .O (syn180329)
    );
    X_BUF \syn20882/XUSED (
      .I (\syn20882/FROM ),
      .O (syn20882)
    );
    defparam C18589.INIT = 16'hFF80;
    X_LUT4 C18589(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [13]),
      .ADR1 (\bridge/configuration/pci_base_addr1 [13]),
      .ADR2 (syn60110),
      .ADR3 (\bridge/configuration/C2001 ),
      .O (\syn180373/GROM )
    );
    defparam C18588.INIT = 16'hFEFC;
    X_LUT4 C18588(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (syn20893),
      .ADR2 (syn180365),
      .ADR3 (\bridge/configuration/pci_err_addr [13]),
      .O (\syn180373/FROM )
    );
    X_BUF \syn180373/YUSED (
      .I (\syn180373/GROM ),
      .O (syn180365)
    );
    X_BUF \syn180373/XUSED (
      .I (\syn180373/FROM ),
      .O (syn180373)
    );
    defparam C18584.INIT = 16'hECA0;
    X_LUT4 C18584(
      .ADR0 (\bridge/configuration/wb_err_addr [13]),
      .ADR1 (\bridge/configuration/C1967 ),
      .ADR2 (\bridge/configuration/C1937 ),
      .ADR3 (\bridge/configuration/pci_err_data [13]),
      .O (\syn180374/GROM )
    );
    defparam C18583.INIT = 16'hFFFE;
    X_LUT4 C18583(
      .ADR0 (syn180366),
      .ADR1 (syn180367),
      .ADR2 (syn180369),
      .ADR3 (syn180368),
      .O (\syn180374/FROM )
    );
    X_BUF \syn180374/YUSED (
      .I (\syn180374/GROM ),
      .O (syn180369)
    );
    X_BUF \syn180374/XUSED (
      .I (\syn180374/FROM ),
      .O (syn180374)
    );
    defparam C18581.INIT = 16'hECA0;
    X_LUT4 C18581(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [13]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_data_out [13]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .O (\syn20922/GROM )
    );
    defparam C18580.INIT = 16'h3230;
    X_LUT4 C18580(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180381),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [13]),
      .O (\syn20922/FROM )
    );
    X_BUF \syn20922/YUSED (
      .I (\syn20922/GROM ),
      .O (syn180381)
    );
    X_BUF \syn20922/XUSED (
      .I (\syn20922/FROM ),
      .O (syn20922)
    );
    defparam C18579.INIT = 16'hC000;
    X_LUT4 C18579(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_base_addr0 [13]),
      .ADR2 (syn16929),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn180387/GROM )
    );
    defparam C18578.INIT = 16'hF8F0;
    X_LUT4 C18578(
      .ADR0 (syn17101),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn20911),
      .ADR3 (\bridge/conf_latency_tim_out [5]),
      .O (\syn180387/FROM )
    );
    X_BUF \syn180387/YUSED (
      .I (\syn180387/GROM ),
      .O (syn20911)
    );
    X_BUF \syn180387/XUSED (
      .I (\syn180387/FROM ),
      .O (syn180387)
    );
    defparam C18572.INIT = 16'hF888;
    X_LUT4 C18572(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [14]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_data_out [14]),
      .ADR3 (syn20493),
      .O (\syn20963/GROM )
    );
    defparam C18571.INIT = 16'h5450;
    X_LUT4 C18571(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [14]),
      .ADR2 (syn180432),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\syn20963/FROM )
    );
    X_BUF \syn20963/YUSED (
      .I (\syn20963/GROM ),
      .O (syn180432)
    );
    X_BUF \syn20963/XUSED (
      .I (\syn20963/FROM ),
      .O (syn20963)
    );
    defparam C18554.INIT = 16'hEAC0;
    X_LUT4 C18554(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [15]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [15]),
      .O (\syn21003/GROM )
    );
    defparam C18553.INIT = 16'h00F8;
    X_LUT4 C18553(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [15]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn180482),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn21003/FROM )
    );
    X_BUF \syn21003/YUSED (
      .I (\syn21003/GROM ),
      .O (syn180482)
    );
    X_BUF \syn21003/XUSED (
      .I (\syn21003/FROM ),
      .O (syn21003)
    );
    defparam C18536.INIT = 16'hFF80;
    X_LUT4 C18536(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [16]),
      .ADR1 (syn60110),
      .ADR2 (\bridge/configuration/pci_base_addr1 [16]),
      .ADR3 (\bridge/configuration/C2001 ),
      .O (\syn180528/GROM )
    );
    defparam C18535.INIT = 16'hFEFC;
    X_LUT4 C18535(
      .ADR0 (\bridge/configuration/pci_err_addr [16]),
      .ADR1 (syn21014),
      .ADR2 (syn180520),
      .ADR3 (\bridge/configuration/C1971 ),
      .O (\syn180528/FROM )
    );
    X_BUF \syn180528/YUSED (
      .I (\syn180528/GROM ),
      .O (syn180520)
    );
    X_BUF \syn180528/XUSED (
      .I (\syn180528/FROM ),
      .O (syn180528)
    );
    defparam C18531.INIT = 16'hECA0;
    X_LUT4 C18531(
      .ADR0 (\bridge/configuration/pci_err_data [16]),
      .ADR1 (\bridge/configuration/wb_err_addr [16]),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (\bridge/configuration/C1937 ),
      .O (\syn180529/GROM )
    );
    defparam C18530.INIT = 16'hFFFE;
    X_LUT4 C18530(
      .ADR0 (syn180523),
      .ADR1 (syn180521),
      .ADR2 (syn180524),
      .ADR3 (syn180522),
      .O (\syn180529/FROM )
    );
    X_BUF \syn180529/YUSED (
      .I (\syn180529/GROM ),
      .O (syn180524)
    );
    X_BUF \syn180529/XUSED (
      .I (\syn180529/FROM ),
      .O (syn180529)
    );
    defparam C18525.INIT = 16'hEAC0;
    X_LUT4 C18525(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [16]),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [16]),
      .O (\syn21041/GROM )
    );
    defparam C18524.INIT = 16'hFCF0;
    X_LUT4 C18524(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [16]),
      .ADR2 (syn180500),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .O (\syn21041/FROM )
    );
    X_BUF \syn21041/YUSED (
      .I (\syn21041/GROM ),
      .O (syn180500)
    );
    X_BUF \syn21041/XUSED (
      .I (\syn21041/FROM ),
      .O (syn21041)
    );
    defparam C18521.INIT = 16'hEAC0;
    X_LUT4 C18521(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [17]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [17]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (syn20493),
      .O (\syn21080/GROM )
    );
    defparam C18520.INIT = 16'h00F8;
    X_LUT4 C18520(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [17]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn180577),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn21080/FROM )
    );
    X_BUF \syn21080/YUSED (
      .I (\syn21080/GROM ),
      .O (syn180577)
    );
    X_BUF \syn21080/XUSED (
      .I (\syn21080/FROM ),
      .O (syn21080)
    );
    defparam C18518.INIT = 16'hFF80;
    X_LUT4 C18518(
      .ADR0 (syn60110),
      .ADR1 (\bridge/configuration/pci_base_addr1 [17]),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [17]),
      .ADR3 (\bridge/configuration/C2001 ),
      .O (\syn180569/GROM )
    );
    defparam C18517.INIT = 16'hFEFA;
    X_LUT4 C18517(
      .ADR0 (syn21053),
      .ADR1 (\bridge/configuration/pci_err_addr [17]),
      .ADR2 (syn180561),
      .ADR3 (\bridge/configuration/C1971 ),
      .O (\syn180569/FROM )
    );
    X_BUF \syn180569/YUSED (
      .I (\syn180569/GROM ),
      .O (syn180561)
    );
    X_BUF \syn180569/XUSED (
      .I (\syn180569/FROM ),
      .O (syn180569)
    );
    defparam C18513.INIT = 16'hF888;
    X_LUT4 C18513(
      .ADR0 (\bridge/configuration/pci_err_data [17]),
      .ADR1 (\bridge/configuration/C1967 ),
      .ADR2 (\bridge/configuration/wb_err_addr [17]),
      .ADR3 (\bridge/configuration/C1937 ),
      .O (\syn180570/GROM )
    );
    defparam C18512.INIT = 16'hFFFE;
    X_LUT4 C18512(
      .ADR0 (syn180562),
      .ADR1 (syn180563),
      .ADR2 (syn180565),
      .ADR3 (syn180564),
      .O (\syn180570/FROM )
    );
    X_BUF \syn180570/YUSED (
      .I (\syn180570/GROM ),
      .O (syn180565)
    );
    X_BUF \syn180570/XUSED (
      .I (\syn180570/FROM ),
      .O (syn180570)
    );
    defparam C18499.INIT = 16'hFFFE;
    X_LUT4 C18499(
      .ADR0 (syn180608),
      .ADR1 (syn180610),
      .ADR2 (syn180611),
      .ADR3 (syn180609),
      .O (\syn21104/GROM )
    );
    defparam C18498.INIT = 16'hFFFE;
    X_LUT4 C18498(
      .ADR0 (syn48754),
      .ADR1 (syn21091),
      .ADR2 (syn180616),
      .ADR3 (syn180607),
      .O (\syn21104/FROM )
    );
    X_BUF \syn21104/YUSED (
      .I (\syn21104/GROM ),
      .O (syn180616)
    );
    X_BUF \syn21104/XUSED (
      .I (\syn21104/FROM ),
      .O (syn21104)
    );
    defparam C18494.INIT = 16'hFF80;
    X_LUT4 C18494(
      .ADR0 (syn16927),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn17063),
      .ADR3 (syn180626),
      .O (\syn180628/GROM )
    );
    defparam C18493.INIT = 16'hF8F0;
    X_LUT4 C18493(
      .ADR0 (\bridge/configuration/pci_base_addr0 [18]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180627),
      .ADR3 (syn16929),
      .O (\syn180628/FROM )
    );
    X_BUF \syn180628/YUSED (
      .I (\syn180628/GROM ),
      .O (syn180627)
    );
    X_BUF \syn180628/XUSED (
      .I (\syn180628/FROM ),
      .O (syn180628)
    );
    defparam C18478.INIT = 16'hF888;
    X_LUT4 C18478(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [19]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (syn20493),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [19]),
      .O (\syn21158/GROM )
    );
    defparam C18477.INIT = 16'hFAF0;
    X_LUT4 C18477(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (VCC),
      .ADR2 (syn180637),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [19]),
      .O (\syn21158/FROM )
    );
    X_BUF \syn21158/YUSED (
      .I (\syn21158/GROM ),
      .O (syn180637)
    );
    X_BUF \syn21158/XUSED (
      .I (\syn21158/FROM ),
      .O (syn21158)
    );
    defparam C18474.INIT = 16'hECA0;
    X_LUT4 C18474(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [20]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_data_out [20]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (syn20493),
      .O (\syn21197/GROM )
    );
    defparam C18473.INIT = 16'h5450;
    X_LUT4 C18473(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn180714),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [20]),
      .O (\syn21197/FROM )
    );
    X_BUF \syn21197/YUSED (
      .I (\syn21197/GROM ),
      .O (syn180714)
    );
    X_BUF \syn21197/XUSED (
      .I (\syn21197/FROM ),
      .O (syn21197)
    );
    defparam C18471.INIT = 16'hFF80;
    X_LUT4 C18471(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [20]),
      .ADR1 (syn60110),
      .ADR2 (\bridge/configuration/pci_base_addr1 [20]),
      .ADR3 (\bridge/configuration/C2001 ),
      .O (\syn180706/GROM )
    );
    defparam C18470.INIT = 16'hFFF8;
    X_LUT4 C18470(
      .ADR0 (\bridge/configuration/pci_err_addr [20]),
      .ADR1 (\bridge/configuration/C1971 ),
      .ADR2 (syn180698),
      .ADR3 (syn21170),
      .O (\syn180706/FROM )
    );
    X_BUF \syn180706/YUSED (
      .I (\syn180706/GROM ),
      .O (syn180698)
    );
    X_BUF \syn180706/XUSED (
      .I (\syn180706/FROM ),
      .O (syn180706)
    );
    defparam C18466.INIT = 16'hF888;
    X_LUT4 C18466(
      .ADR0 (\bridge/configuration/C1937 ),
      .ADR1 (\bridge/configuration/wb_err_addr [20]),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (\bridge/configuration/pci_err_data [20]),
      .O (\syn180707/GROM )
    );
    defparam C18465.INIT = 16'hFFFE;
    X_LUT4 C18465(
      .ADR0 (syn180700),
      .ADR1 (syn180699),
      .ADR2 (syn180702),
      .ADR3 (syn180701),
      .O (\syn180707/FROM )
    );
    X_BUF \syn180707/YUSED (
      .I (\syn180707/GROM ),
      .O (syn180702)
    );
    X_BUF \syn180707/XUSED (
      .I (\syn180707/FROM ),
      .O (syn180707)
    );
    defparam C18458.INIT = 16'hEAC0;
    X_LUT4 C18458(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_data_out [21]),
      .ADR2 (syn20493),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [21]),
      .O (\syn21235/GROM )
    );
    defparam C18457.INIT = 16'h3230;
    X_LUT4 C18457(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180760),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [21]),
      .O (\syn21235/FROM )
    );
    X_BUF \syn21235/YUSED (
      .I (\syn21235/GROM ),
      .O (syn180760)
    );
    X_BUF \syn21235/XUSED (
      .I (\syn21235/FROM ),
      .O (syn21235)
    );
    defparam C18455.INIT = 16'hEAAA;
    X_LUT4 C18455(
      .ADR0 (\bridge/configuration/C2001 ),
      .ADR1 (\bridge/configuration/pci_base_addr1 [21]),
      .ADR2 (syn60110),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [21]),
      .O (\syn180752/GROM )
    );
    defparam C18454.INIT = 16'hFEFA;
    X_LUT4 C18454(
      .ADR0 (syn21208),
      .ADR1 (\bridge/configuration/C1971 ),
      .ADR2 (syn180744),
      .ADR3 (\bridge/configuration/pci_err_addr [21]),
      .O (\syn180752/FROM )
    );
    X_BUF \syn180752/YUSED (
      .I (\syn180752/GROM ),
      .O (syn180744)
    );
    X_BUF \syn180752/XUSED (
      .I (\syn180752/FROM ),
      .O (syn180752)
    );
    defparam C18450.INIT = 16'hEAC0;
    X_LUT4 C18450(
      .ADR0 (\bridge/configuration/wb_err_addr [21]),
      .ADR1 (\bridge/configuration/C1967 ),
      .ADR2 (\bridge/configuration/pci_err_data [21]),
      .ADR3 (\bridge/configuration/C1937 ),
      .O (\syn180753/GROM )
    );
    defparam C18449.INIT = 16'hFFFE;
    X_LUT4 C18449(
      .ADR0 (syn180745),
      .ADR1 (syn180746),
      .ADR2 (syn180748),
      .ADR3 (syn180747),
      .O (\syn180753/FROM )
    );
    X_BUF \syn180753/YUSED (
      .I (\syn180753/GROM ),
      .O (syn180748)
    );
    X_BUF \syn180753/XUSED (
      .I (\syn180753/FROM ),
      .O (syn180753)
    );
    defparam C18436.INIT = 16'hFFFE;
    X_LUT4 C18436(
      .ADR0 (syn180792),
      .ADR1 (syn180793),
      .ADR2 (syn180791),
      .ADR3 (syn180794),
      .O (\syn21259/GROM )
    );
    defparam C18435.INIT = 16'hFFFE;
    X_LUT4 C18435(
      .ADR0 (syn48754),
      .ADR1 (syn21246),
      .ADR2 (syn180799),
      .ADR3 (syn180790),
      .O (\syn21259/FROM )
    );
    X_BUF \syn21259/YUSED (
      .I (\syn21259/GROM ),
      .O (syn180799)
    );
    X_BUF \syn21259/XUSED (
      .I (\syn21259/FROM ),
      .O (syn21259)
    );
    defparam C18431.INIT = 16'hFF80;
    X_LUT4 C18431(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn17059),
      .ADR2 (syn16927),
      .ADR3 (syn180809),
      .O (\syn180811/GROM )
    );
    defparam C18430.INIT = 16'hF8F0;
    X_LUT4 C18430(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn16929),
      .ADR2 (syn180810),
      .ADR3 (\bridge/configuration/pci_base_addr0 [22]),
      .O (\syn180811/FROM )
    );
    X_BUF \syn180811/YUSED (
      .I (\syn180811/GROM ),
      .O (syn180810)
    );
    X_BUF \syn180811/XUSED (
      .I (\syn180811/FROM ),
      .O (syn180811)
    );
    defparam C18415.INIT = 16'hECA0;
    X_LUT4 C18415(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [23]),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [23]),
      .O (\syn21313/GROM )
    );
    defparam C18414.INIT = 16'hFAF0;
    X_LUT4 C18414(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR1 (VCC),
      .ADR2 (syn180820),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [23]),
      .O (\syn21313/FROM )
    );
    X_BUF \syn21313/YUSED (
      .I (\syn21313/GROM ),
      .O (syn180820)
    );
    X_BUF \syn21313/XUSED (
      .I (\syn21313/FROM ),
      .O (syn21313)
    );
    defparam C18404.INIT = 16'hFFFE;
    X_LUT4 C18404(
      .ADR0 (syn180884),
      .ADR1 (syn180885),
      .ADR2 (syn180886),
      .ADR3 (syn180887),
      .O (\syn21346/GROM )
    );
    defparam C18403.INIT = 16'hCCC8;
    X_LUT4 C18403(
      .ADR0 (syn180888),
      .ADR1 (syn181260),
      .ADR2 (syn180892),
      .ADR3 (syn21325),
      .O (\syn21346/FROM )
    );
    X_BUF \syn21346/YUSED (
      .I (\syn21346/GROM ),
      .O (syn180892)
    );
    X_BUF \syn21346/XUSED (
      .I (\syn21346/FROM ),
      .O (syn21346)
    );
    defparam C18410.INIT = 16'hECA0;
    X_LUT4 C18410(
      .ADR0 (\bridge/configuration/C1987 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [24]),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [24]),
      .ADR3 (\bridge/configuration/C1951 ),
      .O (\syn180888/GROM )
    );
    defparam C18409.INIT = 16'hFEFC;
    X_LUT4 C18409(
      .ADR0 (syn60110),
      .ADR1 (\bridge/configuration/C2001 ),
      .ADR2 (syn180883),
      .ADR3 (syn17057),
      .O (\syn180888/FROM )
    );
    X_BUF \syn180888/YUSED (
      .I (\syn180888/GROM ),
      .O (syn180883)
    );
    X_BUF \syn180888/XUSED (
      .I (\syn180888/FROM ),
      .O (syn180888)
    );
    defparam C18400.INIT = 16'h8000;
    X_LUT4 C18400(
      .ADR0 (\bridge/conf_pci_ba1_out [12]),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn16927),
      .ADR3 (\bridge/conf_pci_am1_out [12]),
      .O (\syn180906/GROM )
    );
    defparam C18399.INIT = 16'hF8F0;
    X_LUT4 C18399(
      .ADR0 (\bridge/configuration/status_bit8 ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn21342),
      .ADR3 (syn17098),
      .O (\syn180906/FROM )
    );
    X_BUF \syn180906/YUSED (
      .I (\syn180906/GROM ),
      .O (syn21342)
    );
    X_BUF \syn180906/XUSED (
      .I (\syn180906/FROM ),
      .O (syn180906)
    );
    defparam C18387.INIT = 16'hFFFE;
    X_LUT4 C18387(
      .ADR0 (syn180939),
      .ADR1 (syn180936),
      .ADR2 (syn180937),
      .ADR3 (syn180938),
      .O (\syn21385/GROM )
    );
    defparam C18386.INIT = 16'hCCC8;
    X_LUT4 C18386(
      .ADR0 (syn180940),
      .ADR1 (syn181260),
      .ADR2 (syn180944),
      .ADR3 (syn21365),
      .O (\syn21385/FROM )
    );
    X_BUF \syn21385/YUSED (
      .I (\syn21385/GROM ),
      .O (syn180944)
    );
    X_BUF \syn21385/XUSED (
      .I (\syn21385/FROM ),
      .O (syn21385)
    );
    defparam C18393.INIT = 16'hEAC0;
    X_LUT4 C18393(
      .ADR0 (\bridge/configuration/C1987 ),
      .ADR1 (\bridge/configuration/C1951 ),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [25]),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [25]),
      .O (\syn180940/GROM )
    );
    defparam C18392.INIT = 16'hFFF8;
    X_LUT4 C18392(
      .ADR0 (syn17056),
      .ADR1 (syn60110),
      .ADR2 (syn180935),
      .ADR3 (\bridge/configuration/C2001 ),
      .O (\syn180940/FROM )
    );
    X_BUF \syn180940/YUSED (
      .I (\syn180940/GROM ),
      .O (syn180935)
    );
    X_BUF \syn180940/XUSED (
      .I (\syn180940/FROM ),
      .O (syn180940)
    );
    defparam C18381.INIT = 16'hF800;
    X_LUT4 C18381(
      .ADR0 (syn17056),
      .ADR1 (syn16927),
      .ADR2 (syn17098),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn180961/GROM )
    );
    defparam C18380.INIT = 16'hFFF8;
    X_LUT4 C18380(
      .ADR0 (syn17116),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180958),
      .ADR3 (syn180957),
      .O (\syn180961/FROM )
    );
    X_BUF \syn180961/YUSED (
      .I (\syn180961/GROM ),
      .O (syn180958)
    );
    X_BUF \syn180961/XUSED (
      .I (\syn180961/FROM ),
      .O (syn180961)
    );
    defparam C18353.INIT = 16'hFFEE;
    X_LUT4 C18353(
      .ADR0 (syn181037),
      .ADR1 (syn21448),
      .ADR2 (VCC),
      .ADR3 (syn181038),
      .O (\syn21462/GROM )
    );
    defparam C18352.INIT = 16'hFFFE;
    X_LUT4 C18352(
      .ADR0 (syn181039),
      .ADR1 (syn181040),
      .ADR2 (syn181046),
      .ADR3 (syn181045),
      .O (\syn21462/FROM )
    );
    X_BUF \syn21462/YUSED (
      .I (\syn21462/GROM ),
      .O (syn181046)
    );
    X_BUF \syn21462/XUSED (
      .I (\syn21462/FROM ),
      .O (syn21462)
    );
    defparam C18358.INIT = 16'hECA0;
    X_LUT4 C18358(
      .ADR0 (\bridge/configuration/C1967 ),
      .ADR1 (\bridge/configuration/pci_err_addr [27]),
      .ADR2 (\bridge/configuration/pci_err_data [27]),
      .ADR3 (\bridge/configuration/C1971 ),
      .O (\syn181045/GROM )
    );
    defparam C18357.INIT = 16'hFEFC;
    X_LUT4 C18357(
      .ADR0 (\bridge/configuration/C1973 ),
      .ADR1 (syn48754),
      .ADR2 (syn181041),
      .ADR3 (\bridge/configuration/pci_err_cs_bit31_24 [27]),
      .O (\syn181045/FROM )
    );
    X_BUF \syn181045/YUSED (
      .I (\syn181045/GROM ),
      .O (syn181041)
    );
    X_BUF \syn181045/XUSED (
      .I (\syn181045/FROM ),
      .O (syn181045)
    );
    defparam C18351.INIT = 16'hEAC0;
    X_LUT4 C18351(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [27]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [27]),
      .ADR3 (syn20493),
      .O (\syn21479/GROM )
    );
    defparam C18350.INIT = 16'h5450;
    X_LUT4 C18350(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn181054),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [27]),
      .O (\syn21479/FROM )
    );
    X_BUF \syn21479/YUSED (
      .I (\syn21479/GROM ),
      .O (syn181054)
    );
    X_BUF \syn21479/XUSED (
      .I (\syn21479/FROM ),
      .O (syn21479)
    );
    defparam C18345.INIT = 16'hFF80;
    X_LUT4 C18345(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn16929),
      .ADR2 (\bridge/conf_pci_ba0_out [15]),
      .ADR3 (syn181058),
      .O (\syn181062/GROM )
    );
    defparam C18344.INIT = 16'hFFFE;
    X_LUT4 C18344(
      .ADR0 (syn21465),
      .ADR1 (syn120365),
      .ADR2 (syn181060),
      .ADR3 (syn21466),
      .O (\syn181062/FROM )
    );
    X_BUF \syn181062/YUSED (
      .I (\syn181062/GROM ),
      .O (syn181060)
    );
    X_BUF \syn181062/XUSED (
      .I (\syn181062/FROM ),
      .O (syn181062)
    );
    defparam C18777.INIT = 16'h4040;
    X_LUT4 C18777(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/configuration/C2003 ),
      .ADR2 (syn17106),
      .ADR3 (VCC),
      .O (\syn21465/GROM )
    );
    defparam C18349.INIT = 16'h8080;
    X_LUT4 C18349(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/configuration/status_bit15_11 [11]),
      .ADR2 (syn17098),
      .ADR3 (VCC),
      .O (\syn21465/FROM )
    );
    X_BUF \syn21465/YUSED (
      .I (\syn21465/GROM ),
      .O (syn17098)
    );
    X_BUF \syn21465/XUSED (
      .I (\syn21465/FROM ),
      .O (syn21465)
    );
    defparam C18765.INIT = 16'h0008;
    X_LUT4 C18765(
      .ADR0 (syn16914),
      .ADR1 (\bridge/configuration/C2240 ),
      .ADR2 (\bridge/pciu_conf_offset_out [6]),
      .ADR3 (\bridge/pciu_conf_offset_out [7]),
      .O (\syn120365/GROM )
    );
    defparam C18347.INIT = 16'hC0C0;
    X_LUT4 C18347(
      .ADR0 (VCC),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn17104),
      .ADR3 (VCC),
      .O (\syn120365/FROM )
    );
    X_BUF \syn120365/YUSED (
      .I (\syn120365/GROM ),
      .O (syn17104)
    );
    X_BUF \syn120365/XUSED (
      .I (\syn120365/FROM ),
      .O (syn120365)
    );
    defparam C18334.INIT = 16'hFFFE;
    X_LUT4 C18334(
      .ADR0 (syn181092),
      .ADR1 (syn181094),
      .ADR2 (syn181095),
      .ADR3 (syn181093),
      .O (\syn21511/GROM )
    );
    defparam C18333.INIT = 16'hAAA8;
    X_LUT4 C18333(
      .ADR0 (syn181260),
      .ADR1 (syn181096),
      .ADR2 (syn181100),
      .ADR3 (syn21490),
      .O (\syn21511/FROM )
    );
    X_BUF \syn21511/YUSED (
      .I (\syn21511/GROM ),
      .O (syn181100)
    );
    X_BUF \syn21511/XUSED (
      .I (\syn21511/FROM ),
      .O (syn21511)
    );
    defparam C18340.INIT = 16'hF888;
    X_LUT4 C18340(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [28]),
      .ADR1 (\bridge/configuration/C1951 ),
      .ADR2 (\bridge/configuration/C1987 ),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [28]),
      .O (\syn181096/GROM )
    );
    defparam C18339.INIT = 16'hFFF8;
    X_LUT4 C18339(
      .ADR0 (syn17053),
      .ADR1 (syn60110),
      .ADR2 (syn181091),
      .ADR3 (\bridge/configuration/C2001 ),
      .O (\syn181096/FROM )
    );
    X_BUF \syn181096/YUSED (
      .I (\syn181096/GROM ),
      .O (syn181091)
    );
    X_BUF \syn181096/XUSED (
      .I (\syn181096/FROM ),
      .O (syn181096)
    );
    defparam C18328.INIT = 16'h8080;
    X_LUT4 C18328(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn17098),
      .ADR2 (\bridge/configuration/status_bit15_11 [12]),
      .ADR3 (VCC),
      .O (\syn181114/GROM )
    );
    defparam C18326.INIT = 16'hFEFA;
    X_LUT4 C18326(
      .ADR0 (syn21507),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn21506),
      .ADR3 (syn17104),
      .O (\syn181114/FROM )
    );
    X_BUF \syn181114/YUSED (
      .I (\syn181114/GROM ),
      .O (syn21506)
    );
    X_BUF \syn181114/XUSED (
      .I (\syn181114/FROM ),
      .O (syn181114)
    );
    defparam C18316.INIT = 16'hFFFE;
    X_LUT4 C18316(
      .ADR0 (syn181144),
      .ADR1 (syn181146),
      .ADR2 (syn181145),
      .ADR3 (syn181143),
      .O (\syn21552/GROM )
    );
    defparam C18315.INIT = 16'hAAA8;
    X_LUT4 C18315(
      .ADR0 (syn181260),
      .ADR1 (syn181147),
      .ADR2 (syn181151),
      .ADR3 (syn21531),
      .O (\syn21552/FROM )
    );
    X_BUF \syn21552/YUSED (
      .I (\syn21552/GROM ),
      .O (syn181151)
    );
    X_BUF \syn21552/XUSED (
      .I (\syn21552/FROM ),
      .O (syn21552)
    );
    defparam C18322.INIT = 16'hF888;
    X_LUT4 C18322(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [29]),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [29]),
      .ADR3 (\bridge/configuration/C1987 ),
      .O (\syn181147/GROM )
    );
    defparam C18321.INIT = 16'hFEFA;
    X_LUT4 C18321(
      .ADR0 (\bridge/configuration/C2001 ),
      .ADR1 (syn60110),
      .ADR2 (syn181142),
      .ADR3 (syn17052),
      .O (\syn181147/FROM )
    );
    X_BUF \syn181147/YUSED (
      .I (\syn181147/GROM ),
      .O (syn181142)
    );
    X_BUF \syn181147/XUSED (
      .I (\syn181147/FROM ),
      .O (syn181147)
    );
    defparam C18312.INIT = 16'h8000;
    X_LUT4 C18312(
      .ADR0 (\bridge/conf_pci_ba1_out [17]),
      .ADR1 (syn16927),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (\bridge/conf_pci_am1_out [17]),
      .O (\syn181165/GROM )
    );
    defparam C18311.INIT = 16'hF8F0;
    X_LUT4 C18311(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/configuration/status_bit15_11 [13]),
      .ADR2 (syn21548),
      .ADR3 (syn17098),
      .O (\syn181165/FROM )
    );
    X_BUF \syn181165/YUSED (
      .I (\syn181165/GROM ),
      .O (syn21548)
    );
    X_BUF \syn181165/XUSED (
      .I (\syn181165/FROM ),
      .O (syn181165)
    );
    defparam C18306.INIT = 16'hF888;
    X_LUT4 C18306(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [30]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_data_out [30]),
      .ADR3 (syn20493),
      .O (\syn21601/GROM )
    );
    defparam C18305.INIT = 16'h00F8;
    X_LUT4 C18305(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [30]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn181210),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn21601/FROM )
    );
    X_BUF \syn21601/YUSED (
      .I (\syn21601/GROM ),
      .O (syn181210)
    );
    X_BUF \syn21601/XUSED (
      .I (\syn21601/FROM ),
      .O (syn21601)
    );
    defparam C18288.INIT = 16'hECA0;
    X_LUT4 C18288(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [31]),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [31]),
      .O (\syn21641/GROM )
    );
    defparam C18287.INIT = 16'h00F8;
    X_LUT4 C18287(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [31]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C155 ),
      .ADR2 (syn181265),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn21641/FROM )
    );
    X_BUF \syn21641/YUSED (
      .I (\syn21641/GROM ),
      .O (syn181265)
    );
    X_BUF \syn21641/XUSED (
      .I (\syn21641/FROM ),
      .O (syn21641)
    );
    defparam C18187.INIT = 16'h0303;
    X_LUT4 C18187(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_control_out [1]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_control_out [0]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C749/GROM )
    );
    defparam C18186.INIT = 16'hC444;
    X_LUT4 C18186(
      .ADR0 (\CRT/ssvga_wbm_if/S_41/cell0 ),
      .ADR1 (syn177324),
      .ADR2 (syn181420),
      .ADR3 (syn17678),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C749/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/C749/YUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/C749/GROM ),
      .O (syn181420)
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/C749/XUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/C749/FROM ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C749 )
    );
    defparam C19932.INIT = 16'hC000;
    X_LUT4 C19932(
      .ADR0 (VCC),
      .ADR1 (syn177397),
      .ADR2 (syn177396),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .O (\syn181511/GROM )
    );
    defparam C18145.INIT = 16'h8421;
    X_LUT4 C18145(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [4]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C112 ),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C108 ),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [3]),
      .O (\syn181511/FROM )
    );
    X_BUF \syn181511/YUSED (
      .I (\syn181511/GROM ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C108 )
    );
    X_BUF \syn181511/XUSED (
      .I (\syn181511/FROM ),
      .O (syn181511)
    );
    defparam C18132.INIT = 16'hFF33;
    X_LUT4 C18132(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_first_out ),
      .ADR2 (VCC),
      .ADR3 (syn22083),
      .O (\syn22093/GROM )
    );
    defparam C18131.INIT = 16'h0010;
    X_LUT4 C18131(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_wbr_control_out [0]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (syn22184),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/tabort_ff_in ),
      .O (\syn22093/FROM )
    );
    X_BUF \syn22093/YUSED (
      .I (\syn22093/GROM ),
      .O (syn22184)
    );
    X_BUF \syn22093/XUSED (
      .I (\syn22093/FROM ),
      .O (syn22093)
    );
    defparam C19479.INIT = 16'h0004;
    X_LUT4 C19479(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [0]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [2]),
      .O (\syn22083/GROM )
    );
    defparam C18133.INIT = 16'h7F2A;
    X_LUT4 C18133(
      .ADR0 (\bridge/in_reg_stop_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C248 ),
      .ADR3 (\bridge/in_reg_devsel_out ),
      .O (\syn22083/FROM )
    );
    X_BUF \syn22083/YUSED (
      .I (\syn22083/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C248 )
    );
    X_BUF \syn22083/XUSED (
      .I (\syn22083/FROM ),
      .O (syn22083)
    );
    defparam C18127.INIT = 16'h0011;
    X_LUT4 C18127(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main ),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out ),
      .O (\N12382/GROM )
    );
    defparam C18126.INIT = 16'hF0FC;
    X_LUT4 C18126(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out ),
      .ADR2 (syn22101),
      .ADR3 (syn22096),
      .O (\N12382/FROM )
    );
    X_BUF \N12382/YUSED (
      .I (\N12382/GROM ),
      .O (syn22101)
    );
    X_BUF \N12382/XUSED (
      .I (\N12382/FROM ),
      .O (N12382)
    );
    defparam C17895.INIT = 16'h0005;
    X_LUT4 C17895(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/c_state [0]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/c_state [1]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/c_state [2]),
      .O (\bridge/pci_target_unit/wishbone_master/C81/N3/GROM )
    );
    defparam C17894.INIT = 16'hF0C0;
    X_LUT4 C17894(
      .ADR0 (VCC),
      .ADR1 (syn17011),
      .ADR2 (syn22812),
      .ADR3 (syn17020),
      .O (\bridge/pci_target_unit/wishbone_master/C81/N3/FROM )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/C81/N3/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/C81/N3/GROM ),
      .O (syn22812)
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/C81/N3/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/C81/N3/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C81/N3 )
    );
    defparam C19258.INIT = 16'h1111;
    X_LUT4 C19258(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn17011/GROM )
    );
    defparam C19256.INIT = 16'h00A0;
    X_LUT4 C19256(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_transaction_ready_out ),
      .ADR1 (VCC),
      .ADR2 (syn19577),
      .ADR3 (\bridge/conf_pci_err_pending_out ),
      .O (\syn17011/FROM )
    );
    X_BUF \syn17011/YUSED (
      .I (\syn17011/GROM ),
      .O (syn19577)
    );
    X_BUF \syn17011/XUSED (
      .I (\syn17011/FROM ),
      .O (syn17011)
    );
    defparam C17796.INIT = 16'hAA00;
    X_LUT4 C17796(
      .ADR0 (syn22771),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync_comp_req_pending_out ),
      .O (\N12543/GROM )
    );
    defparam C17794.INIT = 16'hF0F1;
    X_LUT4 C17794(
      .ADR0 (\bridge/pci_target_unit/del_sync/comp_done_reg_main ),
      .ADR1 (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg ),
      .ADR2 (syn23126),
      .ADR3 (\bridge/pciu_pci_drcomp_pending_out ),
      .O (\N12543/FROM )
    );
    X_BUF \N12543/YUSED (
      .I (\N12543/GROM ),
      .O (syn23126)
    );
    X_BUF \N12543/XUSED (
      .I (\N12543/FROM ),
      .O (N12543)
    );
    defparam C19204.INIT = 16'h8880;
    X_LUT4 C19204(
      .ADR0 (syn19708),
      .ADR1 (syn19709),
      .ADR2 (syn179112),
      .ADR3 (syn179113),
      .O (\syn22771/GROM )
    );
    defparam C17907.INIT = 16'hABAA;
    X_LUT4 C17907(
      .ADR0 (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out [1]),
      .ADR1 (\bridge/pci_target_unit/del_sync_bc_out [0]),
      .ADR2 (syn19710),
      .ADR3 (syn17090),
      .O (\syn22771/FROM )
    );
    X_BUF \syn22771/YUSED (
      .I (\syn22771/GROM ),
      .O (syn19710)
    );
    X_BUF \syn22771/XUSED (
      .I (\syn22771/FROM ),
      .O (syn22771)
    );
    defparam C19210.INIT = 16'h003F;
    X_LUT4 C19210(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_burst_out ),
      .ADR2 (\bridge/pci_target_unit/del_sync_bc_out [1]),
      .ADR3 (\bridge/pci_target_unit/del_sync_bc_out [3]),
      .O (\syn19709/GROM )
    );
    defparam C19209.INIT = 16'hFBFF;
    X_LUT4 C19209(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_full_out ),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/almost_full ),
      .ADR2 (syn19701),
      .ADR3 (\bridge/pci_target_unit/del_sync_bc_out [2]),
      .O (\syn19709/FROM )
    );
    X_BUF \syn19709/YUSED (
      .I (\syn19709/GROM ),
      .O (syn19701)
    );
    X_BUF \syn19709/XUSED (
      .I (\syn19709/FROM ),
      .O (syn19709)
    );
    defparam C19208.INIT = 16'h330F;
    X_LUT4 C19208(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync_bc_out [1]),
      .ADR2 (\bridge/pci_target_unit/del_sync_bc_out [3]),
      .ADR3 (\bridge/pci_target_unit/del_sync_burst_out ),
      .O (\syn179112/GROM )
    );
    defparam C19207.INIT = 16'hFFFC;
    X_LUT4 C19207(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/cache_line [6]),
      .ADR2 (syn19698),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/cache_line [5]),
      .O (\syn179112/FROM )
    );
    X_BUF \syn179112/YUSED (
      .I (\syn179112/GROM ),
      .O (syn19698)
    );
    X_BUF \syn179112/XUSED (
      .I (\syn179112/FROM ),
      .O (syn179112)
    );
    defparam C19206.INIT = 16'hFFFE;
    X_LUT4 C19206(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [1]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/cache_line [4]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/cache_line [2]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/cache_line [3]),
      .O (\syn179113/GROM )
    );
    defparam C19205.INIT = 16'hFBFF;
    X_LUT4 C19205(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [7]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/cache_line [0]),
      .ADR2 (syn179111),
      .ADR3 (\bridge/pci_target_unit/del_sync_bc_out [2]),
      .O (\syn179113/FROM )
    );
    X_BUF \syn179113/YUSED (
      .I (\syn179113/GROM ),
      .O (syn179111)
    );
    X_BUF \syn179113/XUSED (
      .I (\syn179113/FROM ),
      .O (syn179113)
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C118 .INIT = 16'hBAAA;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C118 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135 ),
      .ADR1 (N_IRDY),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/N64 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn129 ),
      .O (\bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en/GROM )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C117 .INIT = 16'hFEFA;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C117 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn51 ),
      .ADR1 (N_FRAME),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn137 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/N64 ),
      .O (\bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en/GROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn137 )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/pcit_sm_clk_en )
    );
    defparam C19465.INIT = 16'hFFFE;
    X_LUT4 C19465(
      .ADR0 (syn18899),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C248 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .ADR3 (syn16939),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_sm/state_machine_ce/C42 .INIT = 16'hF4FC;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_sm/state_machine_ce/C42 (
      .ADR0 (N_TRDY),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/ch_state_med ),
      .ADR3 (N_STOP),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/change_state/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/ch_state_med )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/change_state/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state )
    );
    defparam C20011.INIT = 16'h8008;
    X_LUT4 C20011(
      .ADR0 (syn177260),
      .ADR1 (syn176876),
      .ADR2 (\CRT/ssvga_fifo/gray_read_ptr [1]),
      .ADR3 (\CRT/ssvga_fifo/wr_ptr [0]),
      .O (\CRT/ssvga_fifo/S_28/cell0/GROM )
    );
    defparam C20010.INIT = 16'h8000;
    X_LUT4 C20010(
      .ADR0 (syn177262),
      .ADR1 (syn177264),
      .ADR2 (syn177265),
      .ADR3 (syn177263),
      .O (\CRT/ssvga_fifo/S_28/cell0/FROM )
    );
    X_BUF \CRT/ssvga_fifo/S_28/cell0/YUSED (
      .I (\CRT/ssvga_fifo/S_28/cell0/GROM ),
      .O (syn177265)
    );
    X_BUF \CRT/ssvga_fifo/S_28/cell0/XUSED (
      .I (\CRT/ssvga_fifo/S_28/cell0/FROM ),
      .O (\CRT/ssvga_fifo/S_28/cell0 )
    );
    defparam C20019.INIT = 16'h3C3C;
    X_LUT4 C20019(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/gray_read_ptr [6]),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr [4]),
      .ADR3 (VCC),
      .O (\syn177262/GROM )
    );
    defparam C20018.INIT = 16'h6009;
    X_LUT4 C20018(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr [6]),
      .ADR1 (\CRT/ssvga_fifo/gray_read_ptr [7]),
      .ADR2 (syn177249),
      .ADR3 (\CRT/ssvga_fifo/wr_ptr [5]),
      .O (\syn177262/FROM )
    );
    X_BUF \syn177262/YUSED (
      .I (\syn177262/GROM ),
      .O (syn177249)
    );
    X_BUF \syn177262/XUSED (
      .I (\syn177262/FROM ),
      .O (syn177262)
    );
    defparam C20017.INIT = 16'h5A5A;
    X_LUT4 C20017(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr [2]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/gray_read_ptr [4]),
      .ADR3 (VCC),
      .O (\syn177263/GROM )
    );
    defparam C20016.INIT = 16'h4281;
    X_LUT4 C20016(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr [4]),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr [3]),
      .ADR2 (syn177253),
      .ADR3 (\CRT/ssvga_fifo/gray_read_ptr [5]),
      .O (\syn177263/FROM )
    );
    X_BUF \syn177263/YUSED (
      .I (\syn177263/GROM ),
      .O (syn177253)
    );
    X_BUF \syn177263/XUSED (
      .I (\syn177263/FROM ),
      .O (syn177263)
    );
    defparam C20015.INIT = 16'h0FF0;
    X_LUT4 C20015(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/gray_read_ptr [2]),
      .ADR3 (\CRT/ssvga_fifo/wr_ptr [0]),
      .O (\syn177264/GROM )
    );
    defparam C20014.INIT = 16'h4281;
    X_LUT4 C20014(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr [2]),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr [1]),
      .ADR2 (syn177257),
      .ADR3 (\CRT/ssvga_fifo/gray_read_ptr [3]),
      .O (\syn177264/FROM )
    );
    X_BUF \syn177264/YUSED (
      .I (\syn177264/GROM ),
      .O (syn177257)
    );
    X_BUF \syn177264/XUSED (
      .I (\syn177264/FROM ),
      .O (syn177264)
    );
    defparam C20009.INIT = 16'h0002;
    X_LUT4 C20009(
      .ADR0 (\CRT/go ),
      .ADR1 (\CRT/crtc_vblank ),
      .ADR2 (\CRT/ssvga_fifo/S_28/cell0 ),
      .ADR3 (\CRT/crtc_hblank ),
      .O (\CRT/ssvga_fifo/C6/N54/GROM )
    );
    defparam C20008.INIT = 16'hFA0A;
    X_LUT4 C20008(
      .ADR0 (\CRT/ssvga_fifo/rd_ptr [9]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr_plus1 [9]),
      .O (\CRT/ssvga_fifo/C6/N54/FROM )
    );
    X_BUF \CRT/ssvga_fifo/C6/N54/YUSED (
      .I (\CRT/ssvga_fifo/C6/N54/GROM ),
      .O (\CRT/ssvga_fifo/S_45/cell0 )
    );
    X_BUF \CRT/ssvga_fifo/C6/N54/XUSED (
      .I (\CRT/ssvga_fifo/C6/N54/FROM ),
      .O (\CRT/ssvga_fifo/C6/N54 )
    );
    defparam C19937.INIT = 16'h0A00;
    X_LUT4 C19937(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .O (\syn17811/GROM )
    );
    defparam C19933.INIT = 16'h8080;
    X_LUT4 C19933(
      .ADR0 (\bridge/configuration/wb_err_addr [31]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR2 (syn58393),
      .ADR3 (VCC),
      .O (\syn17811/FROM )
    );
    X_BUF \syn17811/YUSED (
      .I (\syn17811/GROM ),
      .O (syn58393)
    );
    X_BUF \syn17811/XUSED (
      .I (\syn17811/FROM ),
      .O (syn17811)
    );
    defparam C19467.INIT = 16'h0020;
    X_LUT4 C19467(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .ADR2 (\bridge/out_bckp_frame_out ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep/GROM )
    );
    defparam C19452.INIT = 16'hF000;
    X_LUT4 C19452(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/frame_en_keep ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_bc_out [0]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/frame_en_keep )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/ad_en_keep )
    );
    defparam C19136.INIT = 16'hAAFF;
    X_LUT4 C19136(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pcit_if_pcir_fifo_data_err_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/devs_w_frm/GROM )
    );
    defparam C19135.INIT = 16'h20A8;
    X_LUT4 C19135(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR2 (syn19959),
      .ADR3 (\bridge/out_bckp_devsel_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/devs_w_frm/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/devs_w_frm/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/devs_w_frm/GROM ),
      .O (syn19959)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/devs_w_frm/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/devs_w_frm/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/devs_w_frm )
    );
    defparam C18890.INIT = 16'h8C84;
    X_LUT4 C18890(
      .ADR0 (\bridge/pciu_conf_offset_out [6]),
      .ADR1 (syn20368),
      .ADR2 (\bridge/pciu_conf_offset_out [5]),
      .ADR3 (\bridge/pciu_conf_offset_out [4]),
      .O (\syn20373/GROM )
    );
    defparam C18889.INIT = 16'hC080;
    X_LUT4 C18889(
      .ADR0 (syn20367),
      .ADR1 (syn20371),
      .ADR2 (syn179679),
      .ADR3 (\bridge/pciu_conf_offset_out [3]),
      .O (\syn20373/FROM )
    );
    X_BUF \syn20373/YUSED (
      .I (\syn20373/GROM ),
      .O (syn179679)
    );
    X_BUF \syn20373/XUSED (
      .I (\syn20373/FROM ),
      .O (syn20373)
    );
    defparam C18731.INIT = 16'h3000;
    X_LUT4 C18731(
      .ADR0 (VCC),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C2240 ),
      .ADR3 (syn60111),
      .O (\syn179986/GROM )
    );
    defparam C18730.INIT = 16'hEAC0;
    X_LUT4 C18730(
      .ADR0 (syn17102),
      .ADR1 (\bridge/configuration/interrupt_line [3]),
      .ADR2 (syn17105),
      .ADR3 (\bridge/conf_cache_line_size_out [3]),
      .O (\syn179986/FROM )
    );
    X_BUF \syn179986/YUSED (
      .I (\syn179986/GROM ),
      .O (syn17105)
    );
    X_BUF \syn179986/XUSED (
      .I (\syn179986/FROM ),
      .O (syn179986)
    );
    defparam C18713.INIT = 16'hB080;
    X_LUT4 C18713(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [4]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR2 (syn19366),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [4]),
      .O (\syn180030/GROM )
    );
    defparam C18712.INIT = 16'hF8F0;
    X_LUT4 C18712(
      .ADR0 (\bridge/configuration/C1929 ),
      .ADR1 (syn16916),
      .ADR2 (syn180029),
      .ADR3 (\bridge/configuration/config_addr[4] ),
      .O (\syn180030/FROM )
    );
    X_BUF \syn180030/YUSED (
      .I (\syn180030/GROM ),
      .O (syn180029)
    );
    X_BUF \syn180030/XUSED (
      .I (\syn180030/FROM ),
      .O (syn180030)
    );
    defparam C18677.INIT = 16'h88C0;
    X_LUT4 C18677(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [7]),
      .ADR1 (syn19366),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [7]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .O (\syn180120/GROM )
    );
    defparam C18676.INIT = 16'hF8F0;
    X_LUT4 C18676(
      .ADR0 (\bridge/configuration/config_addr[7] ),
      .ADR1 (\bridge/configuration/C1929 ),
      .ADR2 (syn180119),
      .ADR3 (syn16916),
      .O (\syn180120/FROM )
    );
    X_BUF \syn180120/YUSED (
      .I (\syn180120/GROM ),
      .O (syn180119)
    );
    X_BUF \syn180120/XUSED (
      .I (\syn180120/FROM ),
      .O (syn180120)
    );
    defparam C18663.INIT = 16'h8000;
    X_LUT4 C18663(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (\bridge/configuration/pci_err_addr [8]),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\syn180180/GROM )
    );
    defparam C18662.INIT = 16'hA8A0;
    X_LUT4 C18662(
      .ADR0 (syn60038),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn180162),
      .ADR3 (syn17105),
      .O (\syn180180/FROM )
    );
    X_BUF \syn180180/YUSED (
      .I (\syn180180/GROM ),
      .O (syn180162)
    );
    X_BUF \syn180180/XUSED (
      .I (\syn180180/FROM ),
      .O (syn180180)
    );
    defparam C18696.INIT = 16'h2000;
    X_LUT4 C18696(
      .ADR0 (syn17005),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (syn60111),
      .ADR3 (syn179659),
      .O (\syn180198/GROM )
    );
    defparam C18638.INIT = 16'hFFF8;
    X_LUT4 C18638(
      .ADR0 (syn17102),
      .ADR1 (\bridge/conf_latency_tim_out [1]),
      .ADR2 (syn17121),
      .ADR3 (\bridge/configuration/wb_err_cs_bit10_8 [9]),
      .O (\syn180198/FROM )
    );
    X_BUF \syn180198/YUSED (
      .I (\syn180198/GROM ),
      .O (syn17121)
    );
    X_BUF \syn180198/XUSED (
      .I (\syn180198/FROM ),
      .O (syn180198)
    );
    defparam C18330.INIT = 16'hF888;
    X_LUT4 C18330(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [28]),
      .ADR1 (syn136384),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [28]),
      .ADR3 (syn136386),
      .O (\syn181113/GROM )
    );
    defparam C18329.INIT = 16'hF8F0;
    X_LUT4 C18329(
      .ADR0 (syn16929),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn181111),
      .ADR3 (\bridge/conf_pci_ba0_out [16]),
      .O (\syn181113/FROM )
    );
    X_BUF \syn181113/YUSED (
      .I (\syn181113/GROM ),
      .O (syn181111)
    );
    X_BUF \syn181113/XUSED (
      .I (\syn181113/FROM ),
      .O (syn181113)
    );
    defparam C18122.INIT = 16'h2000;
    X_LUT4 C18122(
      .ADR0 (syn181563),
      .ADR1 (syn17669),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/img_hit [0]),
      .ADR3 (\CRT/ssvga_wbm_if/S_41/cell0 ),
      .O (\N12383/GROM )
    );
    defparam C18121.INIT = 16'hFAFE;
    X_LUT4 C18121(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg ),
      .ADR2 (N12384),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_clr ),
      .O (\N12383/FROM )
    );
    X_BUF \N12383/YUSED (
      .I (\N12383/GROM ),
      .O (N12384)
    );
    X_BUF \N12383/XUSED (
      .I (\N12383/FROM ),
      .O (N12383)
    );
    defparam C18124.INIT = 16'h0400;
    X_LUT4 C18124(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/map ),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/do_del_request ),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .ADR3 (syn177406),
      .O (\syn181563/GROM )
    );
    defparam C18123.INIT = 16'h80C0;
    X_LUT4 C18123(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out ),
      .ADR1 (syn177324),
      .ADR2 (syn181562),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending ),
      .O (\syn181563/FROM )
    );
    X_BUF \syn181563/YUSED (
      .I (\syn181563/GROM ),
      .O (syn181562)
    );
    X_BUF \syn181563/XUSED (
      .I (\syn181563/FROM ),
      .O (syn181563)
    );
    defparam \bridge/parity_checker/perr_en_crit_gen/C73 .INIT = 16'h5A5A;
    X_LUT4 \bridge/parity_checker/perr_en_crit_gen/C73 (
      .ADR0 (N_PAR),
      .ADR1 (VCC),
      .ADR2 (\bridge/parity_checker/non_critical_par ),
      .ADR3 (VCC),
      .O (\N12033/GROM )
    );
    defparam \bridge/parity_checker/perr_en_crit_gen/C71 .INIT = 16'h1333;
    X_LUT4 \bridge/parity_checker/perr_en_crit_gen/C71 (
      .ADR0 (\bridge/parity_checker/perr_generate ),
      .ADR1 (\bridge/parity_checker/pci_perr_en_reg ),
      .ADR2 (\bridge/parity_checker/perr_en_crit_gen/syn112 ),
      .ADR3 (\bridge/conf_perr_response_out ),
      .O (\N12033/FROM )
    );
    X_BUF \N12033/YUSED (
      .I (\N12033/GROM ),
      .O (\bridge/parity_checker/perr_en_crit_gen/syn112 )
    );
    X_BUF \N12033/XUSED (
      .I (\N12033/FROM ),
      .O (N12033)
    );
    defparam \bridge/parity_checker/C1149 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1149 (
      .ADR0 (\bridge/parity_checker/syn3096 ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .ADR3 (\bridge/parity_checker/syn3164 ),
      .O (\bridge/parity_checker/non_critical_par/GROM )
    );
    defparam \bridge/parity_checker/C1142 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1142 (
      .ADR0 (\bridge/parity_checker/syn3174 ),
      .ADR1 (\bridge/parity_checker/syn3156 ),
      .ADR2 (\bridge/parity_checker/syn3166 ),
      .ADR3 (\bridge/parity_checker/syn3083 ),
      .O (\bridge/parity_checker/non_critical_par/FROM )
    );
    X_BUF \bridge/parity_checker/non_critical_par/YUSED (
      .I (\bridge/parity_checker/non_critical_par/GROM ),
      .O (\bridge/parity_checker/syn3166 )
    );
    X_BUF \bridge/parity_checker/non_critical_par/XUSED (
      .I (\bridge/parity_checker/non_critical_par/FROM ),
      .O (\bridge/parity_checker/non_critical_par )
    );
    defparam \bridge/parity_checker/C1153 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1153 (
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .O (\bridge/parity_checker/syn3156/GROM )
    );
    defparam \bridge/parity_checker/C1152 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1152 (
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .ADR2 (\bridge/parity_checker/syn3155 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .O (\bridge/parity_checker/syn3156/FROM )
    );
    X_BUF \bridge/parity_checker/syn3156/YUSED (
      .I (\bridge/parity_checker/syn3156/GROM ),
      .O (\bridge/parity_checker/syn3155 )
    );
    X_BUF \bridge/parity_checker/syn3156/XUSED (
      .I (\bridge/parity_checker/syn3156/FROM ),
      .O (\bridge/parity_checker/syn3156 )
    );
    defparam C20036.INIT = 16'h4400;
    X_LUT4 C20036(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/c_state [2]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/c_state [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/c_state [0]),
      .O (\syn177213/GROM )
    );
    defparam C20035.INIT = 16'h3350;
    X_LUT4 C20035(
      .ADR0 (\bridge/pci_target_unit/del_sync_be_out [3]),
      .ADR1 (\bridge/pci_target_unit/fifos_pciw_cbe_out [3]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .O (\syn177213/FROM )
    );
    X_BUF \syn177213/YUSED (
      .I (\syn177213/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C960 )
    );
    X_BUF \syn177213/XUSED (
      .I (\syn177213/FROM ),
      .O (syn177213)
    );
    defparam C19893.INIT = 16'h77FF;
    X_LUT4 C19893(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [0]),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .O (\syn18066/GROM )
    );
    defparam C19801.INIT = 16'hF000;
    X_LUT4 C19801(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn17745),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [25]),
      .O (\syn18066/FROM )
    );
    X_BUF \syn18066/YUSED (
      .I (\syn18066/GROM ),
      .O (syn17745)
    );
    X_BUF \syn18066/XUSED (
      .I (\syn18066/FROM ),
      .O (syn18066)
    );
    defparam C19409.INIT = 16'h4050;
    X_LUT4 C19409(
      .ADR0 (syn18863),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (syn19064),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N33/GROM )
    );
    defparam C19408.INIT = 16'hF000;
    X_LUT4 C19408(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_waddr [5]),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N33/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N33/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N33/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/C3/N33/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/C3/N33/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/C3/N33 )
    );
    defparam C19328.INIT = 16'h5050;
    X_LUT4 C19328(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR3 (VCC),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135/GROM )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C119 .INIT = 16'hF8F0;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C119 (
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR1 (N_FRAME),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/N59 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135/FROM )
    );
    X_BUF
     \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135/YUSED (
      .I 
      (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135/GROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/N59 )
    );
    X_BUF
     \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135/XUSED (
      .I 
      (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn135 )
    );
    defparam C19301.INIT = 16'h0300;
    X_LUT4 C19301(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/read_completed_reg ),
      .ADR3 (\bridge/pci_target_unit/del_sync/req_comp_pending ),
      .O (\syn178898/GROM )
    );
    defparam C19300.INIT = 16'hF8F0;
    X_LUT4 C19300(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR1 (syn17000),
      .ADR2 (syn19415),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy ),
      .O (\syn178898/FROM )
    );
    X_BUF \syn178898/YUSED (
      .I (\syn178898/GROM ),
      .O (syn19415)
    );
    X_BUF \syn178898/XUSED (
      .I (\syn178898/FROM ),
      .O (syn178898)
    );
    defparam C19253.INIT = 16'hCEEC;
    X_LUT4 C19253(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C977 ),
      .ADR2 (ACK_I),
      .ADR3 (ERR_I),
      .O (\syn19590/GROM )
    );
    defparam C19252.INIT = 16'hFAF0;
    X_LUT4 C19252(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C983 ),
      .ADR1 (VCC),
      .ADR2 (syn179021),
      .ADR3 (syn17011),
      .O (\syn19590/FROM )
    );
    X_BUF \syn19590/YUSED (
      .I (\syn19590/GROM ),
      .O (syn179021)
    );
    X_BUF \syn19590/XUSED (
      .I (\syn19590/FROM ),
      .O (syn19590)
    );
    defparam C17826.INIT = 16'h0002;
    X_LUT4 C17826(
      .ADR0 (syn17020),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/c_state [1]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/c_state [2]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/c_state [0]),
      .O (\N12510/GROM )
    );
    defparam C17822.INIT = 16'hF2F0;
    X_LUT4 C17822(
      .ADR0 (ACK_I),
      .ADR1 (ERR_I),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .O (\N12510/FROM )
    );
    X_BUF \N12510/YUSED (
      .I (\N12510/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C82/C0 )
    );
    X_BUF \N12510/XUSED (
      .I (\N12510/FROM ),
      .O (N12510)
    );
    defparam C19327.INIT = 16'h000C;
    X_LUT4 C19327(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/previous_frame ),
      .ADR2 (\bridge/out_bckp_frame_en_out ),
      .ADR3 (\bridge/in_reg_frame_out ),
      .O (\syn179261/GROM )
    );
    defparam C19155.INIT = 16'hAABA;
    X_LUT4 C19155(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/N59 ),
      .ADR1 (\bridge/in_reg_irdy_out ),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .ADR3 (\bridge/out_bckp_frame_en_out ),
      .O (\syn179261/FROM )
    );
    X_BUF \syn179261/YUSED (
      .I (\syn179261/GROM ),
      .O (\bridge/pci_target_unit/pcit_sm_addr_phase_out )
    );
    X_BUF \syn179261/XUSED (
      .I (\syn179261/FROM ),
      .O (syn179261)
    );
    defparam C19040.INIT = 16'h0001;
    X_LUT4 C19040(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [13]),
      .ADR1 (\CRT/ssvga_wbm_if/vmaddr_r [12]),
      .ADR2 (\CRT/ssvga_wbm_if/vmaddr_r [11]),
      .ADR3 (\CRT/ssvga_wbm_if/vmaddr_r [10]),
      .O (\syn179382/GROM )
    );
    defparam C19039.INIT = 16'h1000;
    X_LUT4 C19039(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [14]),
      .ADR1 (\CRT/ssvga_wbm_if/vmaddr_r [15]),
      .ADR2 (syn179379),
      .ADR3 (syn179376),
      .O (\syn179382/FROM )
    );
    X_BUF \syn179382/YUSED (
      .I (\syn179382/GROM ),
      .O (syn179379)
    );
    X_BUF \syn179382/XUSED (
      .I (\syn179382/FROM ),
      .O (syn179382)
    );
    defparam C18953.INIT = 16'h0300;
    X_LUT4 C18953(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/vcntr [9]),
      .ADR2 (\CRT/ssvga_crtc/line_end2 ),
      .ADR3 (\CRT/ssvga_crtc/line_end1 ),
      .O (\syn16986/GROM )
    );
    defparam C18951.INIT = 16'hC000;
    X_LUT4 C18951(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/vcntr [4]),
      .ADR2 (syn179548),
      .ADR3 (\CRT/ssvga_crtc/vcntr [1]),
      .O (\syn16986/FROM )
    );
    X_BUF \syn16986/YUSED (
      .I (\syn16986/GROM ),
      .O (syn179548)
    );
    X_BUF \syn16986/XUSED (
      .I (\syn16986/FROM ),
      .O (syn16986)
    );
    defparam C18948.INIT = 16'h7FFF;
    X_LUT4 C18948(
      .ADR0 (\CRT/ssvga_crtc/vcntr [6]),
      .ADR1 (\CRT/ssvga_crtc/vcntr [5]),
      .ADR2 (\CRT/ssvga_crtc/vcntr [8]),
      .ADR3 (\CRT/ssvga_crtc/vcntr [7]),
      .O (\syn179572/GROM )
    );
    defparam C18942.INIT = 16'hFDFF;
    X_LUT4 C18942(
      .ADR0 (\CRT/ssvga_crtc/vcntr [2]),
      .ADR1 (\CRT/ssvga_crtc/vcntr [0]),
      .ADR2 (syn16991),
      .ADR3 (\CRT/ssvga_crtc/vcntr [3]),
      .O (\syn179572/FROM )
    );
    X_BUF \syn179572/YUSED (
      .I (\syn179572/GROM ),
      .O (syn16991)
    );
    X_BUF \syn179572/XUSED (
      .I (\syn179572/FROM ),
      .O (syn179572)
    );
    defparam C18841.INIT = 16'h3020;
    X_LUT4 C18841(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (syn18863),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 ),
      .O (\N12237/GROM )
    );
    defparam C18840.INIT = 16'hA0A0;
    X_LUT4 C18840(
      .ADR0 (\bridge/configuration/wb_error_en ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/S_176/cell0 ),
      .ADR3 (VCC),
      .O (\N12237/FROM )
    );
    X_BUF \N12237/YUSED (
      .I (\N12237/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/S_176/cell0 )
    );
    X_BUF \N12237/XUSED (
      .I (\N12237/FROM ),
      .O (N12237)
    );
    defparam C18834.INIT = 16'h8000;
    X_LUT4 C18834(
      .ADR0 (syn179761),
      .ADR1 (syn16934),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (syn179762),
      .O (\bridge/configuration/C281/N3/GROM )
    );
    defparam C18833.INIT = 16'h00F0;
    X_LUT4 C18833(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn16992),
      .ADR3 (\bridge/in_reg_cbe_out [0]),
      .O (\bridge/configuration/C281/N3/FROM )
    );
    X_BUF \bridge/configuration/C281/N3/YUSED (
      .I (\bridge/configuration/C281/N3/GROM ),
      .O (syn16992)
    );
    X_BUF \bridge/configuration/C281/N3/XUSED (
      .I (\bridge/configuration/C281/N3/FROM ),
      .O (\bridge/configuration/C281/N3 )
    );
    defparam C18665.INIT = 16'hB800;
    X_LUT4 C18665(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [8]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [8]),
      .ADR3 (syn19366),
      .O (\syn180181/GROM )
    );
    defparam C18661.INIT = 16'hC8C0;
    X_LUT4 C18661(
      .ADR0 (syn17121),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn59991),
      .ADR3 (syn17106),
      .O (\syn180181/FROM )
    );
    X_BUF \syn180181/YUSED (
      .I (\syn180181/GROM ),
      .O (syn59991)
    );
    X_BUF \syn180181/XUSED (
      .I (\syn180181/FROM ),
      .O (syn180181)
    );
    defparam C19411.INIT = 16'h00AA;
    X_LUT4 C19411(
      .ADR0 (\bridge/in_reg_devsel_out ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/in_reg_stop_out ),
      .O (\syn181624/GROM )
    );
    defparam C18086.INIT = 16'h000D;
    X_LUT4 C18086(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2 ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_wbr_control_out [0]),
      .O (\syn181624/FROM )
    );
    X_BUF \syn181624/YUSED (
      .I (\syn181624/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 )
    );
    X_BUF \syn181624/XUSED (
      .I (\syn181624/FROM ),
      .O (syn181624)
    );
    defparam C19403.INIT = 16'hF0F2;
    X_LUT4 C19403(
      .ADR0 (syn18908),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last ),
      .ADR2 (syn178714),
      .ADR3 (syn18863),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable/GROM )
    );
    defparam C18078.INIT = 16'hF0A0;
    X_LUT4 C18078(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .ADR1 (VCC),
      .ADR2 (syn19081),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable/FROM )
    );
    X_BUF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable/YUSED (
      .I 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable/GROM ),
      .O (syn19081)
    );
    X_BUF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable/XUSED (
      .I 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable )
    );
    defparam C18068.INIT = 16'h00FC;
    X_LUT4 C18068(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/write_req_int ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_rdy_out ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load/GROM )
    );
    defparam C18067.INIT = 16'h3330;
    X_LUT4 C18067(
      .ADR0 (VCC),
      .ADR1 (N12594),
      .ADR2 (syn22226),
      .ADR3 (syn22225),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/data_be_load/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load/GROM ),
      .O (syn22226)
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/data_be_load/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load )
    );
    defparam C17946.INIT = 16'h8421;
    X_LUT4 C17946(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [25]),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [24]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .O (\syn182015/GROM )
    );
    defparam C17945.INIT = 16'h8000;
    X_LUT4 C17945(
      .ADR0 (syn181990),
      .ADR1 (syn181989),
      .ADR2 (syn181991),
      .ADR3 (syn181988),
      .O (\syn182015/FROM )
    );
    X_BUF \syn182015/YUSED (
      .I (\syn182015/GROM ),
      .O (syn181991)
    );
    X_BUF \syn182015/XUSED (
      .I (\syn182015/FROM ),
      .O (syn182015)
    );
    defparam C17941.INIT = 16'h8241;
    X_LUT4 C17941(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [0]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [1]),
      .O (\syn182018/GROM )
    );
    defparam C17940.INIT = 16'h8000;
    X_LUT4 C17940(
      .ADR0 (syn182001),
      .ADR1 (syn182002),
      .ADR2 (syn182003),
      .ADR3 (syn182000),
      .O (\syn182018/FROM )
    );
    X_BUF \syn182018/YUSED (
      .I (\syn182018/GROM ),
      .O (syn182003)
    );
    X_BUF \syn182018/XUSED (
      .I (\syn182018/FROM ),
      .O (syn182018)
    );
    defparam C17905.INIT = 16'h00FD;
    X_LUT4 C17905(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/almost_empty ),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/stretched_empty ),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/empty ),
      .ADR3 (\bridge/pci_target_unit/fifos_pciw_control_out [0]),
      .O (\syn22805/GROM )
    );
    defparam C17900.INIT = 16'hE0C0;
    X_LUT4 C17900(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C1183 ),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C977 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C723 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .O (\syn22805/FROM )
    );
    X_BUF \syn22805/YUSED (
      .I (\syn22805/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C723 )
    );
    X_BUF \syn22805/XUSED (
      .I (\syn22805/FROM ),
      .O (syn22805)
    );
    defparam C17813.INIT = 16'h0010;
    X_LUT4 C17813(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [0]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [1]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [3]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [2]),
      .O (\syn17006/GROM )
    );
    defparam C17804.INIT = 16'h0003;
    X_LUT4 C17804(
      .ADR0 (VCC),
      .ADR1 (ACK_I),
      .ADR2 (syn23069),
      .ADR3 (ERR_I),
      .O (\syn17006/FROM )
    );
    X_BUF \syn17006/YUSED (
      .I (\syn17006/GROM ),
      .O (syn23069)
    );
    X_BUF \syn17006/XUSED (
      .I (\syn17006/FROM ),
      .O (syn17006)
    );
    defparam C19462.INIT = 16'hFDF0;
    X_LUT4 C19462(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_burst_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/read_bound ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame/GROM )
    );
    defparam C19459.INIT = 16'hFEAA;
    X_LUT4 C19459(
      .ADR0 (syn178588),
      .ADR1 (syn18919),
      .ADR2 (syn178584),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame/GROM ),
      .O (syn178584)
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/slow_frame )
    );
    defparam C19970.INIT = 16'hDD77;
    X_LUT4 C19970(
      .ADR0 (\bridge/conf_wb_am1_out [18]),
      .ADR1 (\bridge/conf_wb_ba1_out [18]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [30]),
      .O (\syn177380/GROM )
    );
    defparam C19969.INIT = 16'h8000;
    X_LUT4 C19969(
      .ADR0 (syn60048),
      .ADR1 (syn60047),
      .ADR2 (syn60049),
      .ADR3 (syn60046),
      .O (\syn177380/FROM )
    );
    X_BUF \syn177380/YUSED (
      .I (\syn177380/GROM ),
      .O (syn60049)
    );
    X_BUF \syn177380/XUSED (
      .I (\syn177380/FROM ),
      .O (syn177380)
    );
    defparam C19306.INIT = 16'h2200;
    X_LUT4 C19306(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/rd_from_fifo ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/cnf_progress ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/same_read_reg ),
      .O (\bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy/GROM )
    );
    defparam C19127.INIT = 16'h0040;
    X_LUT4 C19127(
      .ADR0 (\bridge/out_bckp_trdy_out ),
      .ADR1 (\bridge/out_bckp_trdy_en_out ),
      .ADR2 (syn17000),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy/GROM ),
      .O (syn17000)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/load_med_reg_w_irdy )
    );
    defparam C18958.INIT = 16'h0001;
    X_LUT4 C18958(
      .ADR0 (\CRT/ssvga_crtc/hcntr [4]),
      .ADR1 (\CRT/ssvga_crtc/hcntr [3]),
      .ADR2 (syn48756),
      .ADR3 (\CRT/ssvga_crtc/hcntr [1]),
      .O (\N12151/GROM )
    );
    defparam C18957.INIT = 16'h4010;
    X_LUT4 C18957(
      .ADR0 (\CRT/ssvga_crtc/hcntr [0]),
      .ADR1 (\CRT/ssvga_crtc/hcntr [9]),
      .ADR2 (syn179535),
      .ADR3 (\CRT/ssvga_crtc/hcntr [7]),
      .O (\N12151/FROM )
    );
    X_BUF \N12151/YUSED (
      .I (\N12151/GROM ),
      .O (syn179535)
    );
    X_BUF \N12151/XUSED (
      .I (\N12151/FROM ),
      .O (N12151)
    );
    defparam C18896.INIT = 16'h8000;
    X_LUT4 C18896(
      .ADR0 (syn17005),
      .ADR1 (syn17043),
      .ADR2 (\bridge/pciu_conf_offset_out [5]),
      .ADR3 (\bridge/pciu_conf_offset_out [4]),
      .O (\bridge/configuration/C343/N5/GROM )
    );
    defparam C18828.INIT = 16'h0008;
    X_LUT4 C18828(
      .ADR0 (syn179775),
      .ADR1 (syn179776),
      .ADR2 (\bridge/configuration/C1919 ),
      .ADR3 (\bridge/configuration/C1941 ),
      .O (\bridge/configuration/C343/N5/FROM )
    );
    X_BUF \bridge/configuration/C343/N5/YUSED (
      .I (\bridge/configuration/C343/N5/GROM ),
      .O (\bridge/configuration/C1919 )
    );
    X_BUF \bridge/configuration/C343/N5/XUSED (
      .I (\bridge/configuration/C343/N5/FROM ),
      .O (\bridge/configuration/C343/N5 )
    );
    defparam C18811.INIT = 16'hC0C0;
    X_LUT4 C18811(
      .ADR0 (VCC),
      .ADR1 (syn60090),
      .ADR2 (syn60111),
      .ADR3 (VCC),
      .O (\bridge/configuration/C289/N9/GROM )
    );
    defparam C18810.INIT = 16'h0080;
    X_LUT4 C18810(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR2 (syn17100),
      .ADR3 (\bridge/in_reg_cbe_out [0]),
      .O (\bridge/configuration/C289/N9/FROM )
    );
    X_BUF \bridge/configuration/C289/N9/YUSED (
      .I (\bridge/configuration/C289/N9/GROM ),
      .O (syn17100)
    );
    X_BUF \bridge/configuration/C289/N9/XUSED (
      .I (\bridge/configuration/C289/N9/FROM ),
      .O (\bridge/configuration/C289/N9 )
    );
    defparam C17958.INIT = 16'h8241;
    X_LUT4 C17958(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [16]),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [17]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .O (\syn182016/GROM )
    );
    defparam C17957.INIT = 16'h8000;
    X_LUT4 C17957(
      .ADR0 (syn181994),
      .ADR1 (syn181993),
      .ADR2 (syn181995),
      .ADR3 (syn181992),
      .O (\syn182016/FROM )
    );
    X_BUF \syn182016/YUSED (
      .I (\syn182016/GROM ),
      .O (syn181995)
    );
    X_BUF \syn182016/XUSED (
      .I (\syn182016/FROM ),
      .O (syn182016)
    );
    defparam C17953.INIT = 16'h8421;
    X_LUT4 C17953(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [9]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [9]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [8]),
      .O (\syn182017/GROM )
    );
    defparam C17952.INIT = 16'h8000;
    X_LUT4 C17952(
      .ADR0 (syn181997),
      .ADR1 (syn181998),
      .ADR2 (syn181999),
      .ADR3 (syn181996),
      .O (\syn182017/FROM )
    );
    X_BUF \syn182017/YUSED (
      .I (\syn182017/GROM ),
      .O (syn181999)
    );
    X_BUF \syn182017/XUSED (
      .I (\syn182017/FROM ),
      .O (syn182017)
    );
    defparam C17918.INIT = 16'h0808;
    X_LUT4 C17918(
      .ADR0 (syn182052),
      .ADR1 (syn19366),
      .ADR2 (\bridge/in_reg_irdy_out ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pcir_clear/GROM )
    );
    defparam C17917.INIT = 16'hB333;
    X_LUT4 C17917(
      .ADR0 (\bridge/pci_target_unit/del_sync_comp_flush_out ),
      .ADR1 (N_RST),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/S_198/cell0 ),
      .ADR3 (syn19407),
      .O (\bridge/pci_target_unit/fifos/pcir_clear/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_clear/YUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_clear/GROM ),
      .O (\bridge/pci_target_unit/pci_target_if/S_198/cell0 )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_clear/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_clear/FROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_clear )
    );
    defparam C17825.INIT = 16'h0001;
    X_LUT4 C17825(
      .ADR0 (\bridge/conf_cache_line_size_out [3]),
      .ADR1 (\bridge/conf_cache_line_size_out [6]),
      .ADR2 (\bridge/conf_cache_line_size_out [5]),
      .ADR3 (\bridge/conf_cache_line_size_out [4]),
      .O (\syn23022/GROM )
    );
    defparam C17824.INIT = 16'h0010;
    X_LUT4 C17824(
      .ADR0 (\bridge/conf_cache_line_size_out [2]),
      .ADR1 (\bridge/conf_cache_line_size_out [1]),
      .ADR2 (syn182285),
      .ADR3 (\bridge/conf_cache_line_size_out [7]),
      .O (\syn23022/FROM )
    );
    X_BUF \syn23022/YUSED (
      .I (\syn23022/GROM ),
      .O (syn182285)
    );
    X_BUF \syn23022/XUSED (
      .I (\syn23022/FROM ),
      .O (syn23022)
    );
    defparam C17759.INIT = 16'h8421;
    X_LUT4 C17759(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [1]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [1]),
      .O (\syn182406/GROM )
    );
    defparam C17758.INIT = 16'h8020;
    X_LUT4 C17758(
      .ADR0 (syn182403),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [0]),
      .ADR2 (syn182404),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [0]),
      .O (\syn182406/FROM )
    );
    X_BUF \syn182406/YUSED (
      .I (\syn182406/GROM ),
      .O (syn182404)
    );
    X_BUF \syn182406/XUSED (
      .I (\syn182406/FROM ),
      .O (syn182406)
    );
    defparam C17747.INIT = 16'h8421;
    X_LUT4 C17747(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [1]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [1]),
      .O (\syn23263/GROM )
    );
    defparam C17746.INIT = 16'h8020;
    X_LUT4 C17746(
      .ADR0 (syn182423),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [0]),
      .ADR2 (syn182424),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [0]),
      .O (\syn23263/FROM )
    );
    X_BUF \syn23263/YUSED (
      .I (\syn23263/GROM ),
      .O (syn182424)
    );
    X_BUF \syn23263/XUSED (
      .I (\syn23263/FROM ),
      .O (syn23263)
    );
    defparam C17718.INIT = 16'h8421;
    X_LUT4 C17718(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [1]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [0]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [1]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [0]),
      .O (\syn182488/GROM )
    );
    defparam C17717.INIT = 16'h8080;
    X_LUT4 C17717(
      .ADR0 (syn182484),
      .ADR1 (syn182485),
      .ADR2 (syn182486),
      .ADR3 (VCC),
      .O (\syn182488/FROM )
    );
    X_BUF \syn182488/YUSED (
      .I (\syn182488/GROM ),
      .O (syn182486)
    );
    X_BUF \syn182488/XUSED (
      .I (\syn182488/FROM ),
      .O (syn182488)
    );
    defparam C17687.INIT = 16'h8241;
    X_LUT4 C17687(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [2]),
      .O (\syn182538/GROM )
    );
    defparam C17686.INIT = 16'h8040;
    X_LUT4 C17686(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [0]),
      .ADR1 (syn182535),
      .ADR2 (syn182536),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [0]),
      .O (\syn182538/FROM )
    );
    X_BUF \syn182538/YUSED (
      .I (\syn182538/GROM ),
      .O (syn182536)
    );
    X_BUF \syn182538/XUSED (
      .I (\syn182538/FROM ),
      .O (syn182538)
    );
    defparam C17675.INIT = 16'h8421;
    X_LUT4 C17675(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [1]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0/GROM )
    );
    defparam C17674.INIT = 16'h8040;
    X_LUT4 C17674(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [0]),
      .ADR1 (syn182564),
      .ADR2 (syn182565),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [0]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0/YUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0/GROM ),
      .O (syn182565)
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0/XUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0/FROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/S_82/cell0 )
    );
    defparam C17672.INIT = 16'h8241;
    X_LUT4 C17672(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [2]),
      .O (\syn23568/GROM )
    );
    defparam C17671.INIT = 16'h8020;
    X_LUT4 C17671(
      .ADR0 (syn182555),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [0]),
      .ADR2 (syn182556),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [0]),
      .O (\syn23568/FROM )
    );
    X_BUF \syn23568/YUSED (
      .I (\syn23568/GROM ),
      .O (syn182556)
    );
    X_BUF \syn23568/XUSED (
      .I (\syn23568/FROM ),
      .O (syn23568)
    );
    defparam C17667.INIT = 16'h8241;
    X_LUT4 C17667(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [2]),
      .O (\syn182579/GROM )
    );
    defparam C17666.INIT = 16'h9000;
    X_LUT4 C17666(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [0]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [0]),
      .ADR2 (syn182577),
      .ADR3 (syn182576),
      .O (\syn182579/FROM )
    );
    X_BUF \syn182579/YUSED (
      .I (\syn182579/GROM ),
      .O (syn182577)
    );
    X_BUF \syn182579/XUSED (
      .I (\syn182579/FROM ),
      .O (syn182579)
    );
    defparam C17652.INIT = 16'h8421;
    X_LUT4 C17652(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [1]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [2]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0/GROM )
    );
    defparam C17651.INIT = 16'h8020;
    X_LUT4 C17651(
      .ADR0 (syn182610),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [0]),
      .ADR2 (syn182611),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0/GROM ),
      .O (syn182611)
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0/XUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0/FROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_119/cell0 )
    );
    defparam C17633.INIT = 16'h8241;
    X_LUT4 C17633(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [2]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0/GROM )
    );
    defparam C17632.INIT = 16'h8040;
    X_LUT4 C17632(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [0]),
      .ADR1 (syn182650),
      .ADR2 (syn182651),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0/GROM ),
      .O (syn182651)
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0/XUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0/FROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/S_86/cell0 )
    );
    defparam \bridge/parity_checker/C1135 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1135 (
      .ADR0 (\bridge/out_bckp_ad_out [0]),
      .ADR1 (\bridge/out_bckp_ad_out [1]),
      .ADR2 (\bridge/out_bckp_ad_out [5]),
      .ADR3 (\bridge/out_bckp_ad_out [4]),
      .O (\bridge/parity_checker/data_par/GROM )
    );
    defparam \bridge/parity_checker/C1126 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1126 (
      .ADR0 (\bridge/parity_checker/syn3125 ),
      .ADR1 (\bridge/parity_checker/syn3210 ),
      .ADR2 (\bridge/parity_checker/syn3214 ),
      .ADR3 (\bridge/parity_checker/syn3204 ),
      .O (\bridge/parity_checker/data_par/FROM )
    );
    X_BUF \bridge/parity_checker/data_par/YUSED (
      .I (\bridge/parity_checker/data_par/GROM ),
      .O (\bridge/parity_checker/syn3214 )
    );
    X_BUF \bridge/parity_checker/data_par/XUSED (
      .I (\bridge/parity_checker/data_par/FROM ),
      .O (\bridge/parity_checker/data_par )
    );
    defparam \bridge/parity_checker/C1137 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1137 (
      .ADR0 (\bridge/out_bckp_ad_out [20]),
      .ADR1 (\bridge/out_bckp_ad_out [22]),
      .ADR2 (\bridge/out_bckp_ad_out [19]),
      .ADR3 (\bridge/out_bckp_ad_out [21]),
      .O (\bridge/parity_checker/syn3204/GROM )
    );
    defparam \bridge/parity_checker/C1136 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1136 (
      .ADR0 (\bridge/out_bckp_ad_out [23]),
      .ADR1 (\bridge/out_bckp_ad_out [18]),
      .ADR2 (\bridge/parity_checker/syn3203 ),
      .ADR3 (\bridge/out_bckp_ad_out [17]),
      .O (\bridge/parity_checker/syn3204/FROM )
    );
    X_BUF \bridge/parity_checker/syn3204/YUSED (
      .I (\bridge/parity_checker/syn3204/GROM ),
      .O (\bridge/parity_checker/syn3203 )
    );
    X_BUF \bridge/parity_checker/syn3204/XUSED (
      .I (\bridge/parity_checker/syn3204/FROM ),
      .O (\bridge/parity_checker/syn3204 )
    );
    defparam C19451.INIT = 16'hFDFD;
    X_LUT4 C19451(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [1]),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [0]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/wbs_sm_cbe_out[3]/GROM )
    );
    defparam C19367.INIT = 16'h0F0F;
    X_LUT4 C19367(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (N12360),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/wbs_sm_cbe_out[3]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/wbs_sm_cbe_out<3>/YUSED (
      .I (\bridge/wishbone_slave_unit/wbs_sm_cbe_out[3]/GROM ),
      .O (N12360)
    );
    X_BUF \bridge/wishbone_slave_unit/wbs_sm_cbe_out<3>/XUSED (
      .I (\bridge/wishbone_slave_unit/wbs_sm_cbe_out[3]/FROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_cbe_out [3])
    );
    defparam C19363.INIT = 16'hBFBF;
    X_LUT4 C19363(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_bc_out [2]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_bc_out [1]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_bc_out [3]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_control_out[1]/GROM )
    );
    defparam C19362.INIT = 16'hEAEA;
    X_LUT4 C19362(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 ),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (syn19202),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_control_out[1]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_wbr_control_out<1>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_wbr_control_out[1]/GROM ),
      .O (syn19202)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_wbr_control_out<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_wbr_control_out[1]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_control_out [1])
    );
    defparam C18944.INIT = 16'h0001;
    X_LUT4 C18944(
      .ADR0 (\CRT/ssvga_crtc/hcntr [0]),
      .ADR1 (\CRT/ssvga_crtc/hcntr [2]),
      .ADR2 (\CRT/ssvga_crtc/hcntr [5]),
      .ADR3 (\CRT/ssvga_crtc/hcntr [7]),
      .O (\N12164/GROM )
    );
    defparam C18943.INIT = 16'h0040;
    X_LUT4 C18943(
      .ADR0 (\CRT/ssvga_crtc/hcntr [8]),
      .ADR1 (syn20277),
      .ADR2 (syn179567),
      .ADR3 (\CRT/ssvga_crtc/hcntr [9]),
      .O (\N12164/FROM )
    );
    X_BUF \N12164/YUSED (
      .I (\N12164/GROM ),
      .O (syn179567)
    );
    X_BUF \N12164/XUSED (
      .I (\N12164/FROM ),
      .O (N12164)
    );
    defparam C19458.INIT = 16'hFF88;
    X_LUT4 C19458(
      .ADR0 (\bridge/out_bckp_frame_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2 ),
      .O (\bridge/pci_mux_irdy_in/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_sm/irdy_iob_feed/C42 .INIT = 16'hF4FC;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_sm/irdy_iob_feed/C42 (
      .ADR0 (N_STOP),
      .ADR1 (\bridge/out_bckp_frame_out ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/irdy_slow ),
      .ADR3 (N_TRDY),
      .O (\bridge/pci_mux_irdy_in/FROM )
    );
    X_BUF \bridge/pci_mux_irdy_in/YUSED (
      .I (\bridge/pci_mux_irdy_in/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/irdy_slow )
    );
    X_BUF \bridge/pci_mux_irdy_in/XUSED (
      .I (\bridge/pci_mux_irdy_in/FROM ),
      .O (\bridge/pci_mux_irdy_in )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_burst_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_burst_out/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/burst_out_reg (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/pref_en ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/del_sync_burst_out/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync_burst_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_burst_out/FFY/ASYNC_FF_GSR_OR_104 (
      .I0 (\bridge/wishbone_slave_unit/del_sync_burst_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_burst_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_waddr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [4])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next<4>/FFY/SETOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[4]/FFY/SET )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[4]/FFY/SET ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/trdy_asserted_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/trdy_asserted_reg/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/trdy_asserted_reg_reg (
      .I (\bridge/pci_target_unit/pci_target_if/bckp_trdy_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/trdy_asserted_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/trdy_asserted_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/trdy_asserted_reg/FFY/ASYNC_FF_GSR_OR_105 (
      .I0 (\bridge/pci_target_unit/pci_target_if/trdy_asserted_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/trdy_asserted_reg/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync/req_done_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/req_done_reg/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/req_done_reg_reg (
      .I (\bridge/pci_target_unit/del_sync/req_comp_pending_sample ),
      .CLK (CLK_BUFGPed),
      .CE (N12540),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync/req_done_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/req_done_reg )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/req_done_reg/FFY/ASYNC_FF_GSR_OR_106 (
      .I0 (\bridge/pci_target_unit/del_sync/req_done_reg/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync/req_done_reg/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<12>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[12]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<11> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [11]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N74 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[12]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[11] )
    );
    X_OR2 \bridge/configuration/config_addr<12>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[12]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[12]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N74 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[12]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[12] )
    );
    X_OR2 \bridge/configuration/config_addr<12>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[12]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[12]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<22>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[22]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[22]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[21] )
    );
    X_OR2 \bridge/configuration/config_addr<22>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[22]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[22]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[22]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[22] )
    );
    X_OR2 \bridge/configuration/config_addr<22>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[22]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[22]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<14>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[14]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N74 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[14]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[13] )
    );
    X_OR2 \bridge/configuration/config_addr<14>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[14]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[14]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N74 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[14]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[14] )
    );
    X_OR2 \bridge/configuration/config_addr<14>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[14]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[14]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[23]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[23] )
    );
    X_OR2 \bridge/configuration/config_addr<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[15]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N74 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[15] )
    );
    X_OR2 \bridge/configuration/config_addr<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<16>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[16]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[16]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[16] )
    );
    X_OR2 \bridge/configuration/config_addr<16>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[16]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[16]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<18>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[18]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[18]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[17] )
    );
    X_OR2 \bridge/configuration/config_addr<18>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[18]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[18]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[18]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[18] )
    );
    X_OR2 \bridge/configuration/config_addr<18>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[18]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[18]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_addr_mask1<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_addr_mask1[21]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [20])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [21])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_addr_mask1<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_addr_mask1[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [12])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [13])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<20>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[20]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[20]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[19] )
    );
    X_OR2 \bridge/configuration/config_addr<20>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[20]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[20]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[20]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[20] )
    );
    X_OR2 \bridge/configuration/config_addr<20>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[20]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[20]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pciu_err_bc_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_bc_out[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/bc_register_reg<0> (
      .I (\bridge/pci_target_unit/fifos_pciw_cbe_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .SET (GND),
      .RST (\bridge/pciu_err_bc_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_bc_out [0])
    );
    X_OR2 \bridge/pciu_err_bc_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_bc_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_bc_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/bc_register_reg<1> (
      .I (\bridge/pci_target_unit/fifos_pciw_cbe_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .SET (GND),
      .RST (\bridge/pciu_err_bc_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_bc_out [1])
    );
    X_OR2 \bridge/pciu_err_bc_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_bc_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_bc_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_am1_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_am1_out[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<30> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N3 ),
      .SET (\bridge/conf_pci_am1_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/conf_pci_am1_out [18])
    );
    X_OR2 \bridge/conf_pci_am1_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_am1_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_am1_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<31> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N3 ),
      .SET (\bridge/conf_pci_am1_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/conf_pci_am1_out [19])
    );
    X_OR2 \bridge/conf_pci_am1_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_am1_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_am1_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_addr_mask1<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_addr_mask1[23]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [22])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [23])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_addr_mask1<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_addr_mask1[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [14])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [15])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pciu_err_bc_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_err_bc_out[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/bc_register_reg<2> (
      .I (\bridge/pci_target_unit/fifos_pciw_cbe_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .SET (GND),
      .RST (\bridge/pciu_err_bc_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_bc_out [2])
    );
    X_OR2 \bridge/pciu_err_bc_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_bc_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/bc_register_reg<3> (
      .I (\bridge/pci_target_unit/fifos_pciw_cbe_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .SET (GND),
      .RST (\bridge/pciu_err_bc_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_err_bc_out [3])
    );
    X_OR2 \bridge/pciu_err_bc_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_err_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_err_bc_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_am1_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_am1_out[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<24> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N3 ),
      .SET (\bridge/conf_pci_am1_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/conf_pci_am1_out [12])
    );
    X_OR2 \bridge/conf_pci_am1_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_am1_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_am1_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<25> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N3 ),
      .SET (\bridge/conf_pci_am1_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/conf_pci_am1_out [13])
    );
    X_OR2 \bridge/conf_pci_am1_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_am1_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_am1_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_addr_mask1<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_addr_mask1[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [16])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [17])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_am1_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_am1_out[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<26> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N3 ),
      .SET (\bridge/conf_pci_am1_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/conf_pci_am1_out [14])
    );
    X_OR2 \bridge/conf_pci_am1_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_am1_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_am1_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<27> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N3 ),
      .SET (\bridge/conf_pci_am1_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/conf_pci_am1_out [15])
    );
    X_OR2 \bridge/conf_pci_am1_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_am1_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_am1_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_addr_mask1<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_addr_mask1[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [18])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_addr_mask1[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_addr_mask1 [19])
    );
    X_OR2 \bridge/configuration/pci_addr_mask1<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_addr_mask1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_addr_mask1[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_am1_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_am1_out[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_am1_reg<28> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N3 ),
      .SET (\bridge/conf_pci_am1_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/conf_pci_am1_out [16])
    );
    X_OR2 \bridge/conf_pci_am1_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_am1_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_am1_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_am1_reg<29> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C290/N3 ),
      .SET (\bridge/conf_pci_am1_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/conf_pci_am1_out [17])
    );
    X_OR2 \bridge/conf_pci_am1_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_am1_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_am1_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [0])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<1>/FFY/SETOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFY/SET )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFY/SET ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [1])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<1>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [2])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<3>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [3])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<3>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<5>/F .INIT = 16'h0000;
    X_LUT4 \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<5>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<5>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FROM ),
      .O (GLOBAL_LOGIC0_2)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [4])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<5>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr_reg<5> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [5])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<5>/FFX/SETOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFX/SET )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFX/SET ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr[5]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[4]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_sm_bc0_out/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_sm_bc0_out/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/rw_cbe0_reg (
      .I (\bridge/in_reg_cbe_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_sm_bc0_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_sm_bc0_out )
    );
    X_OR2 \bridge/pci_target_unit/pcit_sm_bc0_out/FFY/ASYNC_FF_GSR_OR_107 (
      .I0 (\bridge/pci_target_unit/pcit_sm_bc0_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_sm_bc0_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<1>/F .INIT = 16'h0000;
    X_LUT4 \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<1>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FROM )
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<1>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/SRNOT )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FROM )
      ,
      .O (GLOBAL_LOGIC0_4)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<3>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17643.INIT = 16'h0FF0;
    X_LUT4 C17643(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [0]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [1]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N360 )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one<0>/BXMUX (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/BXNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/N360 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/BXNOT )
      ,
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17681.INIT = 16'h33CC;
    X_LUT4 C17681(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [0]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N344 )
    );
    X_INV \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one<0>/BXMUX (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [0]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/BXNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/N344 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/BXNOT )
      ,
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17713.INIT = 16'h0FF0;
    X_LUT4 C17713(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [1])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [0])
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N271 )
    );
    defparam C19434.INIT = 16'h8888;
    X_LUT4 C19434(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [1])
      ,
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FROM )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<0>/XUSED (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FROM ),
      .O (syn18979)
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<0>/BXMUX (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [0]),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/BXNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/N271 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [1])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<0>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one_reg<0> (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/BXNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [0])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<0>/FFX/SETOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFX/SET )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFX/SET ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17753.INIT = 16'h33CC;
    X_LUT4 C17753(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [0])
      ,
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [1])
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N326 )
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one<0>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/SRNOT )
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one<0>/BXMUX (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [0]),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/BXNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/N326 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one_reg<0> (
      .I 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/BXNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one[0]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_inTransactionCount<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_inTransactionCount<0>/BYMUX (
      .I (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/BYNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_inTransactionCount_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/in_count_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_inTransactionCount [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_inTransactionCount<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_inTransactionCount[0]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<4>/F .INIT = 16'h0000;
    X_LUT4 \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<4>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<4>/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/FROM ),
      .O (GLOBAL_LOGIC0_5)
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/del_sync/comp_rty_exp_clr/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_rty_exp_clr/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_rty_exp_clr_reg (
      .I (\bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_rty_exp_clr )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR_108 (
      .I0 (\bridge/pci_target_unit/del_sync/comp_rty_exp_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR_109 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/conf_addr_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/conf_addr_out [0])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/conf_addr_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/conf_addr_out [1])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/conf_addr_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/conf_addr_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pciu_conf_offset_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_conf_offset_out[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pciu_conf_offset_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_conf_offset_out [2])
    );
    X_OR2 \bridge/pciu_conf_offset_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_conf_offset_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_conf_offset_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<3> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pciu_conf_offset_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_conf_offset_out [3])
    );
    X_OR2 \bridge/pciu_conf_offset_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_conf_offset_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_conf_offset_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[4]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[4]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr_plus_one [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pciu_conf_offset_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_conf_offset_out[5]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<4> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pciu_conf_offset_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_conf_offset_out [4])
    );
    X_OR2 \bridge/pciu_conf_offset_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_conf_offset_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_conf_offset_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<5> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pciu_conf_offset_out[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_conf_offset_out [5])
    );
    X_OR2 \bridge/pciu_conf_offset_out<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_conf_offset_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_conf_offset_out[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pciu_conf_offset_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/pciu_conf_offset_out[7]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<6> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pciu_conf_offset_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_conf_offset_out [6])
    );
    X_OR2 \bridge/pciu_conf_offset_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_conf_offset_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_conf_offset_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/strd_address_reg<7> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pciu_conf_offset_out[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pciu_conf_offset_out [7])
    );
    X_OR2 \bridge/pciu_conf_offset_out<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pciu_conf_offset_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pciu_conf_offset_out[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_ONE \bridge/configuration/status_bit8/LOGIC_ONE_110 (
      .O (\bridge/configuration/status_bit8/LOGIC_ONE )
    );
    X_FF \bridge/configuration/status_bit8_reg (
      .I (\bridge/configuration/status_bit8/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12313),
      .SET (GND),
      .RST (\bridge/configuration/status_bit8/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/status_bit8 )
    );
    X_OR2 \bridge/configuration/status_bit8/FFY/ASYNC_FF_GSR_OR_111 (
      .I0 (\bridge/configuration/delete_status_bit8 ),
      .I1 (GSR),
      .O (\bridge/configuration/status_bit8/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[4]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr_plus_one [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/raddr[4]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[4]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<3> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[4]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[3] )
    );
    X_OR2 \bridge/configuration/config_addr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[4]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[4]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<4> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[4]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[4] )
    );
    X_OR2 \bridge/configuration/config_addr<4>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[4]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[4]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/previous_frame/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/previous_frame/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/previous_frame_reg (
      .I (\bridge/in_reg_frame_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/pci_target_unit/pci_target_sm/previous_frame/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/pci_target_sm/previous_frame )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/previous_frame/FFY/ASYNC_FF_GSR_OR_112 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/previous_frame/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/previous_frame/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<6>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[6]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<5> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[6]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[5] )
    );
    X_OR2 \bridge/configuration/config_addr<6>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[6]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[6]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<6> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[6]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[6] )
    );
    X_OR2 \bridge/configuration/config_addr<6>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[6]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[6]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[7]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<7> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[7] )
    );
    X_OR2 \bridge/configuration/config_addr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<8>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[8]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<8> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N74 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[8]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[8] )
    );
    X_OR2 \bridge/configuration/config_addr<8>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[8]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[8]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_cs_bit31_24<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_cs_bit31_24[25]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_cs_bit31_24_reg<24> (
      .I (\bridge/pciu_err_bc_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_cs_bit31_24[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_cs_bit31_24 [24])
    );
    X_OR2 \bridge/configuration/pci_err_cs_bit31_24<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_cs_bit31_24[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_cs_bit31_24[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_cs_bit31_24_reg<25> (
      .I (\bridge/pciu_err_bc_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_cs_bit31_24[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_cs_bit31_24 [25])
    );
    X_OR2 \bridge/configuration/pci_err_cs_bit31_24<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_cs_bit31_24[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_cs_bit31_24[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<10>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[10]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<9> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [9]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N74 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[10]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[9] )
    );
    X_OR2 \bridge/configuration/config_addr<10>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[10]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[10]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<10> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [10]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N74 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[10]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[10] )
    );
    X_OR2 \bridge/configuration/config_addr<10>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[10]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[10]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_cs_bit31_24<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_cs_bit31_24[27]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_cs_bit31_24_reg<26> (
      .I (\bridge/pciu_err_bc_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_cs_bit31_24[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_cs_bit31_24 [26])
    );
    X_OR2 \bridge/configuration/pci_err_cs_bit31_24<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_cs_bit31_24[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_cs_bit31_24[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_cs_bit31_24_reg<27> (
      .I (\bridge/pciu_err_bc_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_cs_bit31_24[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_cs_bit31_24 [27])
    );
    X_OR2 \bridge/configuration/pci_err_cs_bit31_24<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_cs_bit31_24[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_cs_bit31_24[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/pci_err_data<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[1]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<0> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [0])
    );
    X_OR2 \bridge/configuration/pci_err_data<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<1> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [1])
    );
    X_OR2 \bridge/configuration/pci_err_data<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/pci_err_data<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[3]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<2> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [2])
    );
    X_OR2 \bridge/configuration/pci_err_data<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<3> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [3])
    );
    X_OR2 \bridge/configuration/pci_err_data<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/pci_err_data<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[5]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<4> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [4]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [4])
    );
    X_OR2 \bridge/configuration/pci_err_data<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<5> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [5]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [5])
    );
    X_OR2 \bridge/configuration/pci_err_data<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_waddr<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[0]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_waddr<0>/BYMUX (
      .I (\bridge/pci_target_unit/fifos/pciw_waddr [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[0]/BYNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_waddr<0>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[0]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/waddr_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_waddr[0]/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_waddr[0]/CENOT ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pciw_waddr[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr [0])
    );
    X_OR2 \bridge/pci_target_unit/fifos/pciw_waddr<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_waddr[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pciw_waddr[0]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[7]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<6> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [6]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [6])
    );
    X_OR2 \bridge/configuration/pci_err_data<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<7> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [7]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [7])
    );
    X_OR2 \bridge/configuration/pci_err_data<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/icr_soft_res/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/icr_soft_res/SRNOT )
    );
    X_FF \bridge/configuration/icr_bit31_reg (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C301/N3 ),
      .SET (GND),
      .RST (\bridge/configuration/icr_soft_res/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/icr_soft_res )
    );
    X_OR2 \bridge/configuration/icr_soft_res/FFY/ASYNC_FF_GSR_OR_113 (
      .I0 (\bridge/configuration/icr_soft_res/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/icr_soft_res/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[9]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<8> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [8]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [8])
    );
    X_OR2 \bridge/configuration/pci_err_data<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<9> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [9]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [9])
    );
    X_OR2 \bridge/configuration/pci_err_data<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[9]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[1]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<0> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [0])
    );
    X_OR2 \bridge/configuration/wb_err_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<1> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [1])
    );
    X_OR2 \bridge/configuration/wb_err_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[3]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<2> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [2])
    );
    X_OR2 \bridge/configuration/wb_err_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<3> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [3])
    );
    X_OR2 \bridge/configuration/wb_err_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_base_addr1<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_base_addr1[13]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N84 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [12])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N84 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [13])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_base_addr1<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_base_addr1[21]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [20])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [21])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[5]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<4> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [4]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [4])
    );
    X_OR2 \bridge/configuration/wb_err_addr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<5> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [5]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [5])
    );
    X_OR2 \bridge/configuration/wb_err_addr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_base_addr1<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_base_addr1[15]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N84 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [14])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N84 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [15])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_ba1_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_ba1_out[19]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<30> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N29 ),
      .SET (GND),
      .RST (\bridge/conf_wb_ba1_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_ba1_out [18])
    );
    X_OR2 \bridge/conf_wb_ba1_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_ba1_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_ba1_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<31> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N29 ),
      .SET (GND),
      .RST (\bridge/conf_wb_ba1_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_ba1_out [19])
    );
    X_OR2 \bridge/conf_wb_ba1_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_ba1_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_ba1_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_base_addr1<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_base_addr1[23]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [22])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [23])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[23]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_io_mux/ad_load_low_gen/C0 .INIT = 16'hFA50;
    X_LUT4 \bridge/pci_io_mux/ad_load_low_gen/C0 (
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_mux_mas_load_in ),
      .ADR3 (\bridge/pci_mux_tar_load_in ),
      .O (\bridge/pci_io_mux/ad_load_ctrl_mhigh/GROM )
    );
    defparam \bridge/pci_io_mux/ad_load_mhigh_gen/C40 .INIT = 16'hF5A0;
    X_LUT4 \bridge/pci_io_mux/ad_load_mhigh_gen/C40 (
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_mux_tar_load_in ),
      .ADR3 (\bridge/pci_mux_mas_load_in ),
      .O (\bridge/pci_io_mux/ad_load_ctrl_mhigh/FROM )
    );
    X_BUF \bridge/pci_io_mux/ad_load_ctrl_mhigh/YUSED (
      .I (\bridge/pci_io_mux/ad_load_ctrl_mhigh/GROM ),
      .O (\bridge/pci_io_mux/ad_load_ctrl_low )
    );
    X_BUF \bridge/pci_io_mux/ad_load_ctrl_mhigh/XUSED (
      .I (\bridge/pci_io_mux/ad_load_ctrl_mhigh/FROM ),
      .O (\bridge/pci_io_mux/ad_load_ctrl_mhigh )
    );
    X_INV \bridge/configuration/wb_err_addr<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[7]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<6> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [6]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [6])
    );
    X_OR2 \bridge/configuration/wb_err_addr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<7> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [7]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [7])
    );
    X_OR2 \bridge/configuration/wb_err_addr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_base_addr1<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_base_addr1[17]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [16])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [17])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_ba1_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_ba1_out[13]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<24> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N29 ),
      .SET (GND),
      .RST (\bridge/conf_wb_ba1_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_ba1_out [12])
    );
    X_OR2 \bridge/conf_wb_ba1_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_ba1_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_ba1_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<25> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N29 ),
      .SET (GND),
      .RST (\bridge/conf_wb_ba1_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_ba1_out [13])
    );
    X_OR2 \bridge/conf_wb_ba1_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_ba1_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_ba1_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/raddr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/wb_err_addr<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[9]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<8> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [8]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [8])
    );
    X_OR2 \bridge/configuration/wb_err_addr<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<9> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [9]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [9])
    );
    X_OR2 \bridge/configuration/wb_err_addr<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[9]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_base_addr1<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_base_addr1[19]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [18])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_base_addr1[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_base_addr1 [19])
    );
    X_OR2 \bridge/configuration/wb_base_addr1<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_base_addr1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_base_addr1[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_ba1_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_ba1_out[15]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<26> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N29 ),
      .SET (GND),
      .RST (\bridge/conf_wb_ba1_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_ba1_out [14])
    );
    X_OR2 \bridge/conf_wb_ba1_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_ba1_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_ba1_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<27> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N29 ),
      .SET (GND),
      .RST (\bridge/conf_wb_ba1_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_ba1_out [15])
    );
    X_OR2 \bridge/conf_wb_ba1_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_ba1_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_ba1_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N94 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [12])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N94 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [13])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[21]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N59 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [20])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N59 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [21])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_io_space_enable_out/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_io_space_enable_out/SRNOT )
    );
    X_FF \bridge/configuration/command_bit2_0_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C281/N3 ),
      .SET (GND),
      .RST (\bridge/conf_io_space_enable_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_io_space_enable_out )
    );
    X_OR2 \bridge/conf_io_space_enable_out/FFY/ASYNC_FF_GSR_OR_114 (
      .I0 (\bridge/conf_io_space_enable_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_io_space_enable_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_ba1_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_ba1_out[17]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<28> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N29 ),
      .SET (GND),
      .RST (\bridge/conf_wb_ba1_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_ba1_out [16])
    );
    X_OR2 \bridge/conf_wb_ba1_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_ba1_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_ba1_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ba1_bit31_12_reg<29> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C294/N29 ),
      .SET (GND),
      .RST (\bridge/conf_wb_ba1_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_ba1_out [17])
    );
    X_OR2 \bridge/conf_wb_ba1_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_ba1_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_ba1_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N94 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [14])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N94 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [15])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[23]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N59 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [22])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N59 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [23])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[31]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<30> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [30])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<31> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [31])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_mem_space_enable_out/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_mem_space_enable_out/SRNOT )
    );
    X_FF \bridge/configuration/command_bit2_0_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C281/N3 ),
      .SET (GND),
      .RST (\bridge/conf_mem_space_enable_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_mem_space_enable_out )
    );
    X_OR2 \bridge/conf_mem_space_enable_out/FFY/ASYNC_FF_GSR_OR_115 (
      .I0 (\bridge/conf_mem_space_enable_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_mem_space_enable_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_master_enable_out/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_master_enable_out/SRNOT )
    );
    X_FF \bridge/configuration/command_bit2_0_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C281/N3 ),
      .SET (GND),
      .RST (\bridge/conf_pci_master_enable_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_master_enable_out )
    );
    X_OR2 \bridge/conf_pci_master_enable_out/FFY/ASYNC_FF_GSR_OR_116 (
      .I0 (\bridge/conf_pci_master_enable_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_master_enable_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N59 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [16])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N59 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [17])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[25]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<24> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [24])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<25> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [25])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N59 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [18])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N59 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [19])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[27]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<26> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [26])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<27> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [27])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_tran_addr1<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_tran_addr1[29]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ta1_reg<28> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [28])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ta1_reg<29> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C291/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_tran_addr1[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_tran_addr1 [29])
    );
    X_OR2 \bridge/configuration/pci_tran_addr1<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_tran_addr1[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_tran_addr1[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_error_en/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_error_en/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_cs_bit0_reg (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C292/N3 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_error_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_error_en )
    );
    X_OR2 \bridge/configuration/pci_error_en/FFY/ASYNC_FF_GSR_OR_117 (
      .I0 (\bridge/configuration/pci_error_en/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_error_en/FFY/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_io_mux/ad_en_mhigh_gen/C0 .INIT = 16'h000F;
    X_LUT4 \bridge/pci_io_mux/ad_en_mhigh_gen/C0 (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_mux_mas_ad_en_in ),
      .ADR3 (\bridge/pci_mux_tar_ad_en_in ),
      .O (\N12330/GROM )
    );
    X_BUF \N12330/YUSED (
      .I (\N12330/GROM ),
      .O (N12330)
    );
    defparam \bridge/parity_checker/C1130 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1130 (
      .ADR0 (\bridge/out_bckp_ad_out [12]),
      .ADR1 (\bridge/out_bckp_ad_out [14]),
      .ADR2 (\bridge/out_bckp_ad_out [11]),
      .ADR3 (\bridge/out_bckp_ad_out [13]),
      .O (\bridge/parity_checker/syn3190/GROM )
    );
    X_BUF \bridge/parity_checker/syn3190/YUSED (
      .I (\bridge/parity_checker/syn3190/GROM ),
      .O (\bridge/parity_checker/syn3190 )
    );
    defparam \bridge/parity_checker/C1131 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1131 (
      .ADR0 (\bridge/out_bckp_ad_out [9]),
      .ADR1 (\bridge/out_bckp_ad_out [8]),
      .ADR2 (\bridge/out_bckp_ad_out [6]),
      .ADR3 (\bridge/out_bckp_ad_out [7]),
      .O (\bridge/parity_checker/syn3189/GROM )
    );
    X_BUF \bridge/parity_checker/syn3189/YUSED (
      .I (\bridge/parity_checker/syn3189/GROM ),
      .O (\bridge/parity_checker/syn3189 )
    );
    defparam \bridge/parity_checker/C1123 .INIT = 16'h4000;
    X_LUT4 \bridge/parity_checker/C1123 (
      .ADR0 (\bridge/in_reg_frame_out ),
      .ADR1 (\bridge/parity_checker/frame_dec2 ),
      .ADR2 (\bridge/conf_serr_enable_out ),
      .ADR3 (\bridge/conf_perr_response_out ),
      .O (\syn18670/GROM )
    );
    defparam C19552.INIT = 16'h4040;
    X_LUT4 C19552(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR1 (\bridge/configuration/C2370 ),
      .ADR2 (\bridge/conf_perr_response_out ),
      .ADR3 (VCC),
      .O (\syn18670/FROM )
    );
    X_BUF \syn18670/YUSED (
      .I (\syn18670/GROM ),
      .O (\bridge/parity_checker/serr_generate )
    );
    X_BUF \syn18670/XUSED (
      .I (\syn18670/FROM ),
      .O (syn18670)
    );
    X_INV \CRT/ssvga_fifo/gray_read_ptr<1>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/gray_read_ptr[1]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<0> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [0]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [0])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<1> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [1]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [1])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[1]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/C1150 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1150 (
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [11]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .O (\syn181997/GROM )
    );
    defparam C17955.INIT = 16'h8241;
    X_LUT4 C17955(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [12]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [13]),
      .O (\syn181997/FROM )
    );
    X_BUF \syn181997/YUSED (
      .I (\syn181997/GROM ),
      .O (\bridge/parity_checker/syn3164 )
    );
    X_BUF \syn181997/XUSED (
      .I (\syn181997/FROM ),
      .O (syn181997)
    );
    defparam \bridge/parity_checker/C1151 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1151 (
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [10]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [9]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[0]/GROM )
    );
    defparam C19329.INIT = 16'hFFF0;
    X_LUT4 C19329(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[0]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<0>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[0]/GROM ),
      .O (\bridge/parity_checker/syn3096 )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<0>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[0]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [0])
    );
    X_INV \CRT/ssvga_fifo/gray_read_ptr<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/gray_read_ptr[3]/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<2> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [2]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [2])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<3> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [3]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [3])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/C1145 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1145 (
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .O (\syn182002/GROM )
    );
    defparam C17942.INIT = 16'h8241;
    X_LUT4 C17942(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [2]),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [3]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .O (\syn182002/FROM )
    );
    X_BUF \syn182002/YUSED (
      .I (\syn182002/GROM ),
      .O (\bridge/parity_checker/syn3172 )
    );
    X_BUF \syn182002/XUSED (
      .I (\syn182002/FROM ),
      .O (syn182002)
    );
    defparam \bridge/parity_checker/C1155 .INIT = 16'hCFFF;
    X_LUT4 \bridge/parity_checker/C1155 (
      .ADR0 (VCC),
      .ADR1 (\bridge/parity_checker/perr_sampled ),
      .ADR2 (\bridge/out_bckp_serr_out ),
      .ADR3 (\bridge/out_bckp_perr_out ),
      .O (\N12313/GROM )
    );
    defparam C18821.INIT = 16'hE000;
    X_LUT4 C18821(
      .ADR0 (\bridge/parity_checker/perr_sampled ),
      .ADR1 (\bridge/parity_checker/pci_perr_en_reg ),
      .ADR2 (\bridge/conf_perr_response_out ),
      .ADR3 (\bridge/parity_checker/master_perr_report ),
      .O (\N12313/FROM )
    );
    X_BUF \N12313/YUSED (
      .I (\N12313/GROM ),
      .O (\bridge/parchk_par_err_detect_out )
    );
    X_BUF \N12313/XUSED (
      .I (\N12313/FROM ),
      .O (N12313)
    );
    defparam \bridge/parity_checker/C1139 .INIT = 16'h2F22;
    X_LUT4 \bridge/parity_checker/C1139 (
      .ADR0 (\bridge/out_bckp_irdy_en_out ),
      .ADR1 (\bridge/in_reg_trdy_out ),
      .ADR2 (\bridge/in_reg_irdy_out ),
      .ADR3 (\bridge/out_bckp_trdy_en_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy/GROM )
    );
    defparam C19302.INIT = 16'h00F0;
    X_LUT4 C19302(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/out_bckp_trdy_en_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy/GROM ),
      .O (\bridge/parity_checker/syn415 )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/tar_load_out_w_irdy )
    );
    defparam \CRT/ssvga_fifo/gray_read_ptr<5>/F .INIT = 16'h0000;
    X_LUT4 \CRT/ssvga_fifo/gray_read_ptr<5>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/gray_read_ptr[5]/FROM )
    );
    X_INV \CRT/ssvga_fifo/gray_read_ptr<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/gray_read_ptr[5]/SRNOT )
    );
    X_BUF \CRT/ssvga_fifo/gray_read_ptr<5>/XUSED (
      .I (\CRT/ssvga_fifo/gray_read_ptr[5]/FROM ),
      .O (GLOBAL_LOGIC0_9)
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<4> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [4]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [4])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<5> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [5]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [5])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pcir_waddr<0>/BYMUX (
      .I (\bridge/pci_target_unit/fifos/pcir_waddr [0]),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[0]/BYNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/waddr_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_waddr[0]/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_waddr[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr [0])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_waddr<0>/FFY/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[0]/FFY/RST )
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_waddr<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_waddr[0]/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[0]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam \CRT/ssvga_fifo/gray_read_ptr<7>/G .INIT = 16'hFFFF;
    X_LUT4 \CRT/ssvga_fifo/gray_read_ptr<7>/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/gray_read_ptr[7]/GROM )
    );
    defparam \CRT/ssvga_fifo/gray_read_ptr<7>/F .INIT = 16'h0000;
    X_LUT4 \CRT/ssvga_fifo/gray_read_ptr<7>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/gray_read_ptr[7]/FROM )
    );
    X_INV \CRT/ssvga_fifo/gray_read_ptr<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/gray_read_ptr[7]/SRNOT )
    );
    X_BUF \CRT/ssvga_fifo/gray_read_ptr<7>/YUSED (
      .I (\CRT/ssvga_fifo/gray_read_ptr[7]/GROM ),
      .O (GLOBAL_LOGIC1)
    );
    X_BUF \CRT/ssvga_fifo/gray_read_ptr<7>/XUSED (
      .I (\CRT/ssvga_fifo/gray_read_ptr[7]/FROM ),
      .O (GLOBAL_LOGIC0_8)
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<6> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [6]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [6])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<7> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [7]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [7])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \CRT/ssvga_fifo/gray_read_ptr<9>/F .INIT = 16'h0000;
    X_LUT4 \CRT/ssvga_fifo/gray_read_ptr<9>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/gray_read_ptr[9]/FROM )
    );
    X_INV \CRT/ssvga_fifo/gray_read_ptr<9>/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/gray_read_ptr[9]/SRNOT )
    );
    X_BUF \CRT/ssvga_fifo/gray_read_ptr<9>/XUSED (
      .I (\CRT/ssvga_fifo/gray_read_ptr[9]/FROM ),
      .O (GLOBAL_LOGIC0_3)
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<8> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [8]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [8])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_fifo/gray_read_ptr_reg<9> (
      .I (\CRT/ssvga_fifo/sync_gray_rd_ptr [9]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/gray_read_ptr[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/gray_read_ptr [9])
    );
    X_OR2 \CRT/ssvga_fifo/gray_read_ptr<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/ssvga_fifo/gray_read_ptr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/gray_read_ptr[9]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_waddr<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/SRNOT )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_waddr<0>/BYMUX (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_waddr [0]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/BYNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/waddr_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr [0])
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbw_waddr<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_waddr[0]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/config_addr<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/config_addr[2]/SRNOT )
    );
    X_FF \bridge/configuration/cnf_addr_bit0_reg (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[2]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[0] )
    );
    X_OR2 \bridge/configuration/config_addr<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[2]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cnf_addr_bit23_2_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C299/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/config_addr[2]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/config_addr[2] )
    );
    X_OR2 \bridge/configuration/config_addr<2>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/config_addr[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/config_addr[2]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_addr_mask1<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_addr_mask1[21]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N64 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [20])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N64 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [21])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_addr_mask1<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_addr_mask1[13]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N89 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [12])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N89 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [13])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_addr_mask1<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_addr_mask1[23]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N64 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [22])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N64 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [23])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_am1_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_am1_out[19]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<30> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N24 ),
      .SET (GND),
      .RST (\bridge/conf_wb_am1_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_am1_out [18])
    );
    X_OR2 \bridge/conf_wb_am1_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_am1_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_am1_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<31> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N24 ),
      .SET (GND),
      .RST (\bridge/conf_wb_am1_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_am1_out [19])
    );
    X_OR2 \bridge/conf_wb_am1_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_am1_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_am1_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_addr_mask1<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_addr_mask1[15]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N89 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [14])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N89 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [15])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[15]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_load_critical/C61 .INIT = 16'hF0F4;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_load_critical/C61 (
      .ADR0 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR1 (\bridge/out_bckp_trdy_en_out ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/N59 ),
      .ADR3 (N_IRDY),
      .O (\syn24519/GROM )
    );
    defparam C19305.INIT = 16'h0030;
    X_LUT4 C19305(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .O (\syn24519/FROM )
    );
    X_BUF \syn24519/YUSED (
      .I (\syn24519/GROM ),
      .O (\bridge/pci_mux_tar_load_in )
    );
    X_BUF \syn24519/XUSED (
      .I (\syn24519/FROM ),
      .O (syn24519)
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/req_done_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/req_done_reg/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/req_done_reg_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample ),
      .CLK (CLK_BUFGPed),
      .CE (N12379),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/req_done_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/req_done_reg )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/req_done_reg/FFY/ASYNC_FF_GSR_OR_118 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/req_done_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/req_done_reg/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_am1_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_am1_out[13]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<24> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N24 ),
      .SET (GND),
      .RST (\bridge/conf_wb_am1_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_am1_out [12])
    );
    X_OR2 \bridge/conf_wb_am1_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_am1_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_am1_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<25> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N24 ),
      .SET (GND),
      .RST (\bridge/conf_wb_am1_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_am1_out [13])
    );
    X_OR2 \bridge/conf_wb_am1_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_am1_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_am1_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_addr_mask1<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_addr_mask1[17]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N64 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [16])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N64 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [17])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_addr_mask1<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_addr_mask1[19]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N64 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [18])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N64 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_addr_mask1[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_addr_mask1 [19])
    );
    X_OR2 \bridge/configuration/wb_addr_mask1<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_addr_mask1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_addr_mask1[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_am1_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_am1_out[15]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<26> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N24 ),
      .SET (GND),
      .RST (\bridge/conf_wb_am1_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_am1_out [14])
    );
    X_OR2 \bridge/conf_wb_am1_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_am1_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_am1_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<27> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N24 ),
      .SET (GND),
      .RST (\bridge/conf_wb_am1_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_am1_out [15])
    );
    X_OR2 \bridge/conf_wb_am1_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_am1_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_am1_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<0> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [0])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<1> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [1])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/delete_wb_err_cs_bit8/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/delete_wb_err_cs_bit8/SRNOT )
    );
    X_FF \bridge/configuration/delete_wb_err_cs_bit8_reg (
      .I (\bridge/configuration/C390/N3 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C346/N5 ),
      .SET (\bridge/configuration/delete_wb_err_cs_bit8/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/configuration/delete_wb_err_cs_bit8 )
    );
    X_OR2 \bridge/configuration/delete_wb_err_cs_bit8/FFY/ASYNC_FF_GSR_OR_119 (
      .I0 (\bridge/configuration/delete_wb_err_cs_bit8/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/delete_wb_err_cs_bit8/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/ssvga_crtc/line_end2/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_crtc/line_end2/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/line_end1_reg (
      .I (crt_hsync),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/line_end2/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/line_end1 )
    );
    X_OR2 \CRT/ssvga_crtc/line_end2/FFY/ASYNC_FF_GSR_OR_120 (
      .I0 (\CRT/ssvga_crtc/line_end2/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/line_end2/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_crtc/line_end2_reg (
      .I (\CRT/ssvga_crtc/line_end1 ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_crtc/line_end2/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_crtc/line_end2 )
    );
    X_OR2 \CRT/ssvga_crtc/line_end2/FFX/ASYNC_FF_GSR_OR_121 (
      .I0 (\CRT/ssvga_crtc/line_end2/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_crtc/line_end2/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_am1_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_am1_out[17]/SRNOT )
    );
    X_FF \bridge/configuration/wb_am1_reg<28> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N24 ),
      .SET (GND),
      .RST (\bridge/conf_wb_am1_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_am1_out [16])
    );
    X_OR2 \bridge/conf_wb_am1_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_am1_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_am1_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_am1_reg<29> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C296/N24 ),
      .SET (GND),
      .RST (\bridge/conf_wb_am1_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_am1_out [17])
    );
    X_OR2 \bridge/conf_wb_am1_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_am1_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_am1_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<2> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [2])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<3> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [3])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<4> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [4])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<5> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [5])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[5]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/wb_err_data<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[11]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<10> (
      .I (\bridge/out_bckp_ad_out [10]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [10])
    );
    X_OR2 \bridge/configuration/wb_err_data<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<11> (
      .I (\bridge/out_bckp_ad_out [11]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [11])
    );
    X_OR2 \bridge/configuration/wb_err_data<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[11]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<6> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [6]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [6])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<7> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [7]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [7])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[7]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/wb_err_data<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[21]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<20> (
      .I (\bridge/out_bckp_ad_out [20]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [20])
    );
    X_OR2 \bridge/configuration/wb_err_data<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<21> (
      .I (\bridge/out_bckp_ad_out [21]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [21])
    );
    X_OR2 \bridge/configuration/wb_err_data<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[13]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<12> (
      .I (\bridge/out_bckp_ad_out [12]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [12])
    );
    X_OR2 \bridge/configuration/wb_err_data<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<13> (
      .I (\bridge/out_bckp_ad_out [13]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [13])
    );
    X_OR2 \bridge/configuration/wb_err_data<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<8> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [8]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [8])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<9> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [9]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [9])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[9]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/wb_err_data<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[31]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<30> (
      .I (\bridge/out_bckp_ad_out [30]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [30])
    );
    X_OR2 \bridge/configuration/wb_err_data<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<31> (
      .I (\bridge/out_bckp_ad_out [31]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [31])
    );
    X_OR2 \bridge/configuration/wb_err_data<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[23]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<22> (
      .I (\bridge/out_bckp_ad_out [22]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [22])
    );
    X_OR2 \bridge/configuration/wb_err_data<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<23> (
      .I (\bridge/out_bckp_ad_out [23]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [23])
    );
    X_OR2 \bridge/configuration/wb_err_data<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[15]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<14> (
      .I (\bridge/out_bckp_ad_out [14]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [14])
    );
    X_OR2 \bridge/configuration/wb_err_data<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<15> (
      .I (\bridge/out_bckp_ad_out [15]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [15])
    );
    X_OR2 \bridge/configuration/wb_err_data<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[25]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<24> (
      .I (\bridge/out_bckp_ad_out [24]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [24])
    );
    X_OR2 \bridge/configuration/wb_err_data<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<25> (
      .I (\bridge/out_bckp_ad_out [25]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [25])
    );
    X_OR2 \bridge/configuration/wb_err_data<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[17]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<16> (
      .I (\bridge/out_bckp_ad_out [16]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [16])
    );
    X_OR2 \bridge/configuration/wb_err_data<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<17> (
      .I (\bridge/out_bckp_ad_out [17]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [17])
    );
    X_OR2 \bridge/configuration/wb_err_data<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[27]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<26> (
      .I (\bridge/out_bckp_ad_out [26]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [26])
    );
    X_OR2 \bridge/configuration/wb_err_data<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<27> (
      .I (\bridge/out_bckp_ad_out [27]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [27])
    );
    X_OR2 \bridge/configuration/wb_err_data<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[19]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<18> (
      .I (\bridge/out_bckp_ad_out [18]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [18])
    );
    X_OR2 \bridge/configuration/wb_err_data<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<19> (
      .I (\bridge/out_bckp_ad_out [19]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [19])
    );
    X_OR2 \bridge/configuration/wb_err_data<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[29]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<28> (
      .I (\bridge/out_bckp_ad_out [28]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [28])
    );
    X_OR2 \bridge/configuration/wb_err_data<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<29> (
      .I (\bridge/out_bckp_ad_out [29]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [29])
    );
    X_OR2 \bridge/configuration/wb_err_data<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<0> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [0])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<1> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [1])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<2> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [2])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<3> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [3])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[5]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<4> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [4]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [4])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<5> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [5]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [5])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \crt_hsync/SRMUX (
      .I (N_RST),
      .O (\crt_hsync/SRNOT )
    );
    X_INV \crt_hsync/BYMUX (
      .I (\CRT/ssvga_crtc/hcntr [6]),
      .O (\crt_hsync/BYNOT )
    );
    X_FF \CRT/ssvga_crtc/hsync_reg (
      .I (\crt_hsync/BYNOT ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12164),
      .SET (GND),
      .RST (\crt_hsync/FFY/ASYNC_FF_GSR_OR ),
      .O (crt_hsync)
    );
    X_OR2 \crt_hsync/FFY/ASYNC_FF_GSR_OR_122 (
      .I0 (\crt_hsync/SRNOT ),
      .I1 (GSR),
      .O (\crt_hsync/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<1>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/CENOT ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[7]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<6> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [6]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [6])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<7> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [7]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [7])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<3>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/conf_pci_img_ctrl1_out<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_img_ctrl1_out[0]/SRNOT )
    );
    X_FF \bridge/configuration/pci_img_ctrl1_bit2_1_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C289/N9 ),
      .SET (GND),
      .RST (\bridge/conf_pci_img_ctrl1_out[0]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_img_ctrl1_out [0])
    );
    X_OR2 \bridge/conf_pci_img_ctrl1_out<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_img_ctrl1_out[0]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_img_ctrl1_out[0]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[9]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<8> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [8]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [8])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<9> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [9]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [9])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[9]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_img_ctrl1<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_img_ctrl1[2]/SRNOT )
    );
    X_FF \bridge/configuration/pci_img_ctrl1_bit2_1_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C289/N9 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_img_ctrl1[2]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_img_ctrl1 [2])
    );
    X_OR2 \bridge/configuration/pci_img_ctrl1<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_img_ctrl1[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_img_ctrl1[2]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<4>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/CENOT ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_ONE \bridge/conf_pci_err_pending_out/LOGIC_ONE_123 (
      .O (\bridge/conf_pci_err_pending_out/LOGIC_ONE )
    );
    X_FF \bridge/configuration/pci_err_cs_bit8_reg (
      .I (\bridge/conf_pci_err_pending_out/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/conf_pci_err_pending_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_err_pending_out )
    );
    X_OR2 \bridge/conf_pci_err_pending_out/FFY/ASYNC_FF_GSR_OR_124 (
      .I0 (\bridge/configuration/delete_pci_err_cs_bit8 ),
      .I1 (GSR),
      .O (\bridge/conf_pci_err_pending_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_mem_io1_out/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_mem_io1_out/SRNOT )
    );
    X_FF \bridge/configuration/wb_ba1_bit0_reg (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C295/N3 ),
      .SET (GND),
      .RST (\bridge/conf_wb_mem_io1_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_mem_io1_out )
    );
    X_OR2 \bridge/conf_wb_mem_io1_out/FFY/ASYNC_FF_GSR_OR_125 (
      .I0 (\bridge/conf_wb_mem_io1_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_mem_io1_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[4]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/wishbone_slave_unit/del_sync_bc_out<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/SRNOT )
    );
    X_ONE \bridge/wishbone_slave_unit/del_sync_bc_out<2>/LOGIC_ONE (
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/LOGIC_ONE )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_bc_out<2>/BXMUX (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/map ),
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/BXNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/bc_out_reg<1> (
      .I (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out [1])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_bc_out<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/bc_out_reg<2> (
      .I (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/BXNOT ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/FFX/ASYNC_FF_GSR_OR )
      ,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out [2])
    );
    X_OR2 \bridge/wishbone_slave_unit/del_sync_bc_out<2>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/del_sync_bc_out[2]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_sm/frame_iob_ce/C42 .INIT = 16'hBAFA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_sm/frame_iob_ce/C42 (
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/frame_load_slow ),
      .ADR1 (N_TRDY),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (N_STOP),
      .O (\bridge/wishbone_slave_unit/pcim_sm_first_out/GROM )
    );
    defparam C18227.INIT = 16'hA0A2;
    X_LUT4 C18227(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (N_DEVSEL),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_first_out ),
      .ADR3 (N_TRDY),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/transfer_input )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_sm_first_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_sm_first_out/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_first_out/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_first_out/GROM ),
      .O (\bridge/pci_mux_frame_load_in )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/transfer_reg (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/transfer_input ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/pcim_sm_first_out/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_first_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_sm_first_out/FFX/ASYNC_FF_GSR_OR_126 (
      .I0 (\bridge/wishbone_slave_unit/pcim_sm_first_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_sm_first_out/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<4>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_waddr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/CENOT ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<1>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/CENOT ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/CENOT ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<3>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/CENOT ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<4>/CEMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/CENOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/CENOT ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/pci_err_data<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[11]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<10> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [10]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [10])
    );
    X_OR2 \bridge/configuration/pci_err_data<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<11> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [11]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [11])
    );
    X_OR2 \bridge/configuration/pci_err_data<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[11]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync/sync_comp_done/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/sync_comp_done/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/done_sync/sync_data_out_reg<0> (
      .I (\bridge/pci_target_unit/del_sync/req_done_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/sync_comp_done/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/sync_comp_done )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/sync_comp_done/FFY/ASYNC_FF_GSR_OR_127 (
      .I0 (\bridge/pci_target_unit/del_sync/sync_comp_done/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync/sync_comp_done/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/sync_comp_done/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/sync_comp_done/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/done_sync/sync_data_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/del_sync/req_done_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/sync_comp_done/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/sync_comp_done )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/sync_comp_done/FFY/ASYNC_FF_GSR_OR_128 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/sync_comp_done/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/sync_comp_done/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_bc_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_bc_out[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/bc_out_reg<0> (
      .I (\bridge/pci_target_unit/pcit_if_bc_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_bc_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_bc_out [0])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_bc_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_bc_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_bc_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/bc_out_reg<1> (
      .I (\bridge/pci_target_unit/pcit_if_bc_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_bc_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_bc_out [1])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_bc_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_bc_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_bc_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[21]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<20> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [20]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [20])
    );
    X_OR2 \bridge/configuration/pci_err_data<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<21> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [21]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [21])
    );
    X_OR2 \bridge/configuration/pci_err_data<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<12> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [12]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [12])
    );
    X_OR2 \bridge/configuration/pci_err_data<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<13> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [13]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [13])
    );
    X_OR2 \bridge/configuration/pci_err_data<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_bc_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_bc_out[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/bc_out_reg<2> (
      .I (\bridge/pci_target_unit/pcit_if_bc_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (\bridge/pci_target_unit/del_sync_bc_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/del_sync_bc_out [2])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_bc_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_bc_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/bc_out_reg<3> (
      .I (\bridge/pci_target_unit/pcit_if_bc_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_bc_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_bc_out [3])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_bc_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_bc_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[31]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<30> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [30]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [30])
    );
    X_OR2 \bridge/configuration/pci_err_data<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<31> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [31]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [31])
    );
    X_OR2 \bridge/configuration/pci_err_data<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[23]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<22> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [22]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [22])
    );
    X_OR2 \bridge/configuration/pci_err_data<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<23> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [23]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [23])
    );
    X_OR2 \bridge/configuration/pci_err_data<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<14> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [14]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [14])
    );
    X_OR2 \bridge/configuration/pci_err_data<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<15> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [15]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [15])
    );
    X_OR2 \bridge/configuration/pci_err_data<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_wbr_be_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/SRNOT )
    );
    X_ONE \bridge/wishbone_slave_unit/pcim_if_wbr_be_out<1>/LOGIC_ONE (
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/LOGIC_ONE )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/be_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_wbr_be_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/be_out_reg<1> (
      .I (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_wbr_be_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[25]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<24> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [24]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [24])
    );
    X_OR2 \bridge/configuration/pci_err_data<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<25> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [25]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [25])
    );
    X_OR2 \bridge/configuration/pci_err_data<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<16> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [16]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [16])
    );
    X_OR2 \bridge/configuration/pci_err_data<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<17> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [17]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [17])
    );
    X_OR2 \bridge/configuration/pci_err_data<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_wbr_be_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/SRNOT )
    );
    X_ONE \bridge/wishbone_slave_unit/pcim_if_wbr_be_out<3>/LOGIC_ONE (
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/LOGIC_ONE )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/be_out_reg<2> (
      .I (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_wbr_be_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/be_out_reg<3> (
      .I (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12384),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pcim_if_wbr_be_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pcim_if_wbr_be_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[27]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<26> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [26]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [26])
    );
    X_OR2 \bridge/configuration/pci_err_data<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<27> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [27]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [27])
    );
    X_OR2 \bridge/configuration/pci_err_data<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_data<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<18> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [18]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [18])
    );
    X_OR2 \bridge/configuration/pci_err_data<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<19> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [19]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [19])
    );
    X_OR2 \bridge/configuration/pci_err_data<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/SRNOT )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<0>/BYMUX (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [0]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/BYNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/in_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_inTransactionCount[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/pci_err_data<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_data[29]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_data_reg<28> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [28]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [28])
    );
    X_OR2 \bridge/configuration/pci_err_data<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_data_reg<29> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [29]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_data[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_data [29])
    );
    X_OR2 \bridge/configuration/pci_err_data<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_data[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_data[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \N_LED/SRMUX (
      .I (N_RST),
      .O (\N_LED/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/ctrl_r_reg<0> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12118),
      .SET (GND),
      .RST (\N_LED/FFY/ASYNC_FF_GSR_OR ),
      .O (N_LED)
    );
    X_OR2 \N_LED/FFY/ASYNC_FF_GSR_OR_129 (
      .I0 (\N_LED/SRNOT ),
      .I1 (GSR),
      .O (\N_LED/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[11]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<10> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [10]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [10])
    );
    X_OR2 \bridge/configuration/wb_err_addr<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<11> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [11]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [11])
    );
    X_OR2 \bridge/configuration/wb_err_addr<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[11]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[21]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<20> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [20]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [20])
    );
    X_OR2 \bridge/configuration/wb_err_addr<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<21> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [21]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [21])
    );
    X_OR2 \bridge/configuration/wb_err_addr<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[13]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<12> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [12]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [12])
    );
    X_OR2 \bridge/configuration/wb_err_addr<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<13> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [13]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [13])
    );
    X_OR2 \bridge/configuration/wb_err_addr<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_cs_bit31_24<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_cs_bit31_24[31]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_cs_bit31_24_reg<30> (
      .I (\bridge/out_bckp_cbe_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit31_24[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit31_24 [30])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit31_24<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit31_24[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit31_24[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_cs_bit31_24_reg<31> (
      .I (\bridge/out_bckp_cbe_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit31_24[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit31_24 [31])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit31_24<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit31_24[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit31_24[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[31]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<30> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [30]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [30])
    );
    X_OR2 \bridge/configuration/wb_err_addr<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<31> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [31]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [31])
    );
    X_OR2 \bridge/configuration/wb_err_addr<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[23]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<22> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [22]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [22])
    );
    X_OR2 \bridge/configuration/wb_err_addr<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<23> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [23]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [23])
    );
    X_OR2 \bridge/configuration/wb_err_addr<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[15]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<14> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [14]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [14])
    );
    X_OR2 \bridge/configuration/wb_err_addr<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<15> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [15]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [15])
    );
    X_OR2 \bridge/configuration/wb_err_addr<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_cs_bit31_24<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_cs_bit31_24[25]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_cs_bit31_24_reg<24> (
      .I (\bridge/wishbone_slave_unit/pcim_if_bc_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit31_24[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit31_24 [24])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit31_24<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit31_24[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit31_24[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_cs_bit31_24_reg<25> (
      .I (\bridge/wishbone_slave_unit/pcim_if_bc_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit31_24[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit31_24 [25])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit31_24<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit31_24[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit31_24[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[25]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<24> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [24]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [24])
    );
    X_OR2 \bridge/configuration/wb_err_addr<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<25> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [25]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [25])
    );
    X_OR2 \bridge/configuration/wb_err_addr<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[17]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<16> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [16]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [16])
    );
    X_OR2 \bridge/configuration/wb_err_addr<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<17> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [17]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [17])
    );
    X_OR2 \bridge/configuration/wb_err_addr<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_cs_bit31_24<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_cs_bit31_24[27]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_cs_bit31_24_reg<26> (
      .I (\bridge/wishbone_slave_unit/pcim_if_bc_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit31_24[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit31_24 [26])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit31_24<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit31_24[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit31_24[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_cs_bit31_24_reg<27> (
      .I (\bridge/wishbone_slave_unit/pcim_if_bc_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit31_24[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit31_24 [27])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit31_24<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit31_24[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit31_24[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[27]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<26> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [26]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [26])
    );
    X_OR2 \bridge/configuration/wb_err_addr<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<27> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [27]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [27])
    );
    X_OR2 \bridge/configuration/wb_err_addr<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[19]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<18> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [18]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [18])
    );
    X_OR2 \bridge/configuration/wb_err_addr<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<19> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [19]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [19])
    );
    X_OR2 \bridge/configuration/wb_err_addr<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/ssvga_fifo/rd_ssvga_en/SRMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/rd_ssvga_en/SRNOT )
    );
    X_FF \CRT/ssvga_fifo/rd_ssvga_en_reg (
      .I (\CRT/ssvga_fifo/sync_ssvga_en ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CRT/ssvga_fifo/rd_ssvga_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/ssvga_fifo/rd_ssvga_en )
    );
    X_OR2 \CRT/ssvga_fifo/rd_ssvga_en/FFY/ASYNC_FF_GSR_OR_130 (
      .I0 (\CRT/ssvga_fifo/rd_ssvga_en/SRNOT ),
      .I1 (GSR),
      .O (\CRT/ssvga_fifo/rd_ssvga_en/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_cs_bit31_24<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_cs_bit31_24[29]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_cs_bit31_24_reg<28> (
      .I (\bridge/out_bckp_cbe_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit31_24[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit31_24 [28])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit31_24<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit31_24[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit31_24[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_cs_bit31_24_reg<29> (
      .I (\bridge/out_bckp_cbe_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_cs_bit31_24[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_cs_bit31_24 [29])
    );
    X_OR2 \bridge/configuration/wb_err_cs_bit31_24<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_cs_bit31_24[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_cs_bit31_24[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_addr<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_addr[29]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<28> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [28]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [28])
    );
    X_OR2 \bridge/configuration/wb_err_addr<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_addr_reg<29> (
      .I (\bridge/wishbone_slave_unit/pcim_if_address_out [29]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_addr[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_addr [29])
    );
    X_OR2 \bridge/configuration/wb_err_addr<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_addr[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_addr[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[13]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N84 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [12])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N84 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [13])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[21]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [20])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [21])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/del_sync_be_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_be_out[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/be_out_reg<0> (
      .I (\bridge/in_reg_cbe_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_be_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_be_out [0])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_be_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_be_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_be_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/be_out_reg<1> (
      .I (\bridge/in_reg_cbe_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_be_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_be_out [1])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_be_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_be_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_be_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[15]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N84 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [14])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N84 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [15])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[31]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<30> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [30])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<31> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [31])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[23]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [22])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [23])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/del_sync_be_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_be_out[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/be_out_reg<2> (
      .I (\bridge/in_reg_cbe_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_be_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_be_out [2])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_be_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_be_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_be_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/be_out_reg<3> (
      .I (\bridge/in_reg_cbe_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_be_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_be_out [3])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_be_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_be_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_be_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[17]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [16])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [17])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[25]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<24> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [24])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<25> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [25])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[25]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_io_mux/ad_load_mlow_gen/C0 .INIT = 16'hD8D8;
    X_LUT4 \bridge/pci_io_mux/ad_load_mlow_gen/C0 (
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/pci_mux_tar_load_in ),
      .ADR2 (\bridge/pci_mux_mas_load_in ),
      .ADR3 (VCC),
      .O (\bridge/pci_io_mux/ad_load_ctrl_high/GROM )
    );
    defparam \bridge/pci_io_mux/ad_load_high_gen/C0 .INIT = 16'hCFC0;
    X_LUT4 \bridge/pci_io_mux/ad_load_high_gen/C0 (
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_mux_tar_load_in ),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (\bridge/pci_mux_mas_load_in ),
      .O (\bridge/pci_io_mux/ad_load_ctrl_high/FROM )
    );
    X_BUF \bridge/pci_io_mux/ad_load_ctrl_high/YUSED (
      .I (\bridge/pci_io_mux/ad_load_ctrl_high/GROM ),
      .O (\bridge/pci_io_mux/ad_load_ctrl_mlow )
    );
    X_BUF \bridge/pci_io_mux/ad_load_ctrl_high/XUSED (
      .I (\bridge/pci_io_mux/ad_load_ctrl_high/FROM ),
      .O (\bridge/pci_io_mux/ad_load_ctrl_high )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[4]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus1 [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/wb_tran_addr1<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[27]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<26> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [26])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<27> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [27])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[19]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [18])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N69 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [19])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync/sync_req_rty_exp/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/sync_req_rty_exp/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/rty_exp_sync/sync_data_out_reg<0> (
      .I (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/sync_req_rty_exp/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/sync_req_rty_exp )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/sync_req_rty_exp/FFY/ASYNC_FF_GSR_OR_131 (
      .I0 (\bridge/pci_target_unit/del_sync/sync_req_rty_exp/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/sync_req_rty_exp/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_tran_addr1<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_tran_addr1[29]/SRNOT )
    );
    X_FF \bridge/configuration/wb_ta1_reg<28> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [28])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_ta1_reg<29> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C297/N29 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_tran_addr1[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_tran_addr1 [29])
    );
    X_OR2 \bridge/configuration/wb_tran_addr1<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_tran_addr1[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_tran_addr1[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/crtc_hblank/SRMUX (
      .I (N_RST),
      .O (\CRT/crtc_hblank/SRNOT )
    );
    X_FF \CRT/ssvga_crtc/hblank_reg (
      .I (\CRT/ssvga_crtc/hcntr [9]),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12151),
      .SET (GND),
      .RST (\CRT/crtc_hblank/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/crtc_hblank )
    );
    X_OR2 \CRT/crtc_hblank/FFY/ASYNC_FF_GSR_OR_132 (
      .I0 (\CRT/crtc_hblank/SRNOT ),
      .I1 (GSR),
      .O (\CRT/crtc_hblank/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[1]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr/SRNOT )
    );
    X_FF
     \bridge/pci_target_unit/del_sync/rty_exp_back_prop_sync/sync_data_out_reg<0> (
      .I (\bridge/pci_target_unit/del_sync/req_rty_exp_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR_133 (
      .I0 (\bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/sync_comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/del_sync/rty_exp_back_prop_sync/sync_data_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR_134 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/sync_comp_rty_exp_clr/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus1 [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg_reg<0> (
      .I (\bridge/pci_target_unit/fifos_pcir_control_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg [0])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg_reg<1> (
      .I (\bridge/pci_target_unit/fifos_pcir_control_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg [1])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_ctrl_reg[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \CRT/pix_start_addr<3>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[3]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<2> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [2])
    );
    X_OR2 \CRT/pix_start_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<3> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [3])
    );
    X_OR2 \CRT/pix_start_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[3]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<5>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[5]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<4> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [4]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [4])
    );
    X_OR2 \CRT/pix_start_addr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<5> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [5]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [5])
    );
    X_OR2 \CRT/pix_start_addr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[5]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/parity_checker/master_perr_report/SRMUX (
      .I (N_RST),
      .O (\bridge/parity_checker/master_perr_report/SRNOT )
    );
    X_FF \bridge/parity_checker/master_perr_report_reg (
      .I (\bridge/out_bckp_irdy_en_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/parity_checker/master_perr_report/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/parity_checker/master_perr_report )
    );
    X_OR2 \bridge/parity_checker/master_perr_report/FFY/ASYNC_FF_GSR_OR_135 (
      .I0 (\bridge/parity_checker/master_perr_report/SRNOT ),
      .I1 (GSR),
      .O (\bridge/parity_checker/master_perr_report/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_img_ctrl1<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_img_ctrl1[2]/SRNOT )
    );
    X_FF \bridge/configuration/wb_img_ctrl1_bit2_0_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C293/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_img_ctrl1[2]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_img_ctrl1[0] )
    );
    X_OR2 \bridge/configuration/wb_img_ctrl1<2>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_img_ctrl1[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_img_ctrl1[2]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_img_ctrl1_bit2_0_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C293/N14 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_img_ctrl1[2]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_img_ctrl1[2] )
    );
    X_OR2 \bridge/configuration/wb_img_ctrl1<2>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_img_ctrl1[2]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_img_ctrl1[2]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<7>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[7]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<6> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [6]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [6])
    );
    X_OR2 \CRT/pix_start_addr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<7> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [7]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [7])
    );
    X_OR2 \CRT/pix_start_addr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[7]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_wb_img_ctrl1_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_wb_img_ctrl1_out[1]/SRNOT )
    );
    X_FF \bridge/configuration/wb_img_ctrl1_bit2_0_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C293/N14 ),
      .SET (GND),
      .RST (\bridge/conf_wb_img_ctrl1_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_img_ctrl1_out [1])
    );
    X_OR2 \bridge/conf_wb_img_ctrl1_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_wb_img_ctrl1_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_wb_img_ctrl1_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<9>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[9]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<8> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [8]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [8])
    );
    X_OR2 \CRT/pix_start_addr<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<9> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [9]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [9])
    );
    X_OR2 \CRT/pix_start_addr<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[9]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[9]/FFX/ASYNC_FF_GSR_OR )
    );
    X_ONE \bridge/configuration/status_bit15_11<15>/LOGIC_ONE (
      .O (\bridge/configuration/status_bit15_11[15]/LOGIC_ONE )
    );
    X_FF \bridge/configuration/status_bit15_11_reg<15> (
      .I (\bridge/configuration/status_bit15_11[15]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/parchk_par_err_detect_out ),
      .SET (GND),
      .RST (\bridge/configuration/status_bit15_11[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/status_bit15_11 [15])
    );
    X_OR2 \bridge/configuration/status_bit15_11<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/delete_status_bit15 ),
      .I1 (GSR),
      .O (\bridge/configuration/status_bit15_11[15]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C20001.INIT = 16'hDD88;
    X_LUT4 C20001(
      .ADR0 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [2]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [2]),
      .O (\CRT/ssvga_fifo/C6/N18/GROM )
    );
    defparam C20002.INIT = 16'hD8D8;
    X_LUT4 C20002(
      .ADR0 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [3]),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [3]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C6/N18/FROM )
    );
    X_BUF \CRT/ssvga_fifo/C6/N18/YUSED (
      .I (\CRT/ssvga_fifo/C6/N18/GROM ),
      .O (\CRT/ssvga_fifo/C6/N12 )
    );
    X_BUF \CRT/ssvga_fifo/C6/N18/XUSED (
      .I (\CRT/ssvga_fifo/C6/N18/FROM ),
      .O (\CRT/ssvga_fifo/C6/N18 )
    );
    defparam C20003.INIT = 16'hF0CC;
    X_LUT4 C20003(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr [4]),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr_plus1 [4]),
      .ADR3 (\CRT/ssvga_fifo/S_45/cell0 ),
      .O (\CRT/ssvga_fifo/C6/N30/GROM )
    );
    defparam C20004.INIT = 16'hFA50;
    X_LUT4 C20004(
      .ADR0 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [5]),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr_plus1 [5]),
      .O (\CRT/ssvga_fifo/C6/N30/FROM )
    );
    X_BUF \CRT/ssvga_fifo/C6/N30/YUSED (
      .I (\CRT/ssvga_fifo/C6/N30/GROM ),
      .O (\CRT/ssvga_fifo/C6/N24 )
    );
    X_BUF \CRT/ssvga_fifo/C6/N30/XUSED (
      .I (\CRT/ssvga_fifo/C6/N30/FROM ),
      .O (\CRT/ssvga_fifo/C6/N30 )
    );
    defparam C20021.INIT = 16'hFC0C;
    X_LUT4 C20021(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/dat_o_low [0]),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [1]),
      .ADR3 (\CRT/ssvga_fifo/dat_o_high [0]),
      .O (\CRT/fifo_out[1]/GROM )
    );
    defparam C20022.INIT = 16'hB8B8;
    X_LUT4 C20022(
      .ADR0 (\CRT/ssvga_fifo/dat_o_high [1]),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr [1]),
      .ADR2 (\CRT/ssvga_fifo/dat_o_low [1]),
      .ADR3 (VCC),
      .O (\CRT/fifo_out[1]/FROM )
    );
    X_BUF \CRT/fifo_out<1>/YUSED (
      .I (\CRT/fifo_out[1]/GROM ),
      .O (\CRT/fifo_out [0])
    );
    X_BUF \CRT/fifo_out<1>/XUSED (
      .I (\CRT/fifo_out[1]/FROM ),
      .O (\CRT/fifo_out [1])
    );
    defparam C20013.INIT = 16'h5AA5;
    X_LUT4 C20013(
      .ADR0 (\CRT/ssvga_fifo/gray_read_ptr [8]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr [7]),
      .ADR3 (\CRT/ssvga_fifo/wr_ptr [6]),
      .O (\syn176876/GROM )
    );
    X_BUF \syn176876/YUSED (
      .I (\syn176876/GROM ),
      .O (syn176876)
    );
    defparam C20005.INIT = 16'hDD88;
    X_LUT4 C20005(
      .ADR0 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [6]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [6]),
      .O (\CRT/ssvga_fifo/C6/N42/GROM )
    );
    defparam C20006.INIT = 16'hE4E4;
    X_LUT4 C20006(
      .ADR0 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr [7]),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr_plus1 [7]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/C6/N42/FROM )
    );
    X_BUF \CRT/ssvga_fifo/C6/N42/YUSED (
      .I (\CRT/ssvga_fifo/C6/N42/GROM ),
      .O (\CRT/ssvga_fifo/C6/N36 )
    );
    X_BUF \CRT/ssvga_fifo/C6/N42/XUSED (
      .I (\CRT/ssvga_fifo/C6/N42/FROM ),
      .O (\CRT/ssvga_fifo/C6/N42 )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [0])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<1>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [1])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<1>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[11]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<10> (
      .I (ADR_O[10]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [10])
    );
    X_OR2 \bridge/configuration/pci_err_addr<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<11> (
      .I (\bridge/pciu_err_addr_out[11] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [11])
    );
    X_OR2 \bridge/configuration/pci_err_addr<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C20023.INIT = 16'hAFA0;
    X_LUT4 C20023(
      .ADR0 (\CRT/ssvga_fifo/dat_o_high [2]),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [1]),
      .ADR3 (\CRT/ssvga_fifo/dat_o_low [2]),
      .O (\CRT/fifo_out[3]/GROM )
    );
    defparam C20024.INIT = 16'hCCAA;
    X_LUT4 C20024(
      .ADR0 (\CRT/ssvga_fifo/dat_o_low [3]),
      .ADR1 (\CRT/ssvga_fifo/dat_o_high [3]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [1]),
      .O (\CRT/fifo_out[3]/FROM )
    );
    X_BUF \CRT/fifo_out<3>/YUSED (
      .I (\CRT/fifo_out[3]/GROM ),
      .O (\CRT/fifo_out [2])
    );
    X_BUF \CRT/fifo_out<3>/XUSED (
      .I (\CRT/fifo_out[3]/FROM ),
      .O (\CRT/fifo_out [3])
    );
    defparam C20025.INIT = 16'hCCF0;
    X_LUT4 C20025(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/dat_o_high [4]),
      .ADR2 (\CRT/ssvga_fifo/dat_o_low [4]),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [1]),
      .O (\CRT/fifo_out[5]/GROM )
    );
    defparam C20026.INIT = 16'hCFC0;
    X_LUT4 C20026(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/dat_o_high [5]),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr [1]),
      .ADR3 (\CRT/ssvga_fifo/dat_o_low [5]),
      .O (\CRT/fifo_out[5]/FROM )
    );
    X_BUF \CRT/fifo_out<5>/YUSED (
      .I (\CRT/fifo_out[5]/GROM ),
      .O (\CRT/fifo_out [4])
    );
    X_BUF \CRT/fifo_out<5>/XUSED (
      .I (\CRT/fifo_out[5]/FROM ),
      .O (\CRT/fifo_out [5])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [2])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<3>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [3])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<3>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_sm_rdy_out/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_sm_rdy_out/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/bckp_trdy_reg_reg (
      .I (\bridge/out_bckp_trdy_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\bridge/pci_target_unit/pcit_sm_rdy_out/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/pci_target_unit/pcit_sm_rdy_out )
    );
    X_OR2 \bridge/pci_target_unit/pcit_sm_rdy_out/FFY/ASYNC_FF_GSR_OR_136 (
      .I0 (\bridge/pci_target_unit/pcit_sm_rdy_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_sm_rdy_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[21]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<20> (
      .I (\bridge/pciu_err_addr_out[20] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [20])
    );
    X_OR2 \bridge/configuration/pci_err_addr<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<21> (
      .I (\bridge/pciu_err_addr_out[21] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [21])
    );
    X_OR2 \bridge/configuration/pci_err_addr<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<12> (
      .I (\bridge/pciu_err_addr_out[12] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [12])
    );
    X_OR2 \bridge/configuration/pci_err_addr<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<13> (
      .I (\bridge/pciu_err_addr_out[13] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [13])
    );
    X_OR2 \bridge/configuration/pci_err_addr<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[13]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C20027.INIT = 16'hFC30;
    X_LUT4 C20027(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr [1]),
      .ADR2 (\CRT/ssvga_fifo/dat_o_low [6]),
      .ADR3 (\CRT/ssvga_fifo/dat_o_high [6]),
      .O (\CRT/fifo_out[7]/GROM )
    );
    defparam C20028.INIT = 16'hAACC;
    X_LUT4 C20028(
      .ADR0 (\CRT/ssvga_fifo/dat_o_high [7]),
      .ADR1 (\CRT/ssvga_fifo/dat_o_low [7]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [1]),
      .O (\CRT/fifo_out[7]/FROM )
    );
    X_BUF \CRT/fifo_out<7>/YUSED (
      .I (\CRT/fifo_out[7]/GROM ),
      .O (\CRT/fifo_out [6])
    );
    X_BUF \CRT/fifo_out<7>/XUSED (
      .I (\CRT/fifo_out[7]/FROM ),
      .O (\CRT/fifo_out [7])
    );
    X_INV \bridge/configuration/interrupt_line<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/interrupt_line[1]/SRNOT )
    );
    X_FF \bridge/configuration/interrupt_line_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C288/N39 ),
      .SET (GND),
      .RST (\bridge/configuration/interrupt_line[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/interrupt_line [0])
    );
    X_OR2 \bridge/configuration/interrupt_line<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/interrupt_line[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/interrupt_line[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/interrupt_line_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C288/N39 ),
      .SET (GND),
      .RST (\bridge/configuration/interrupt_line[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/interrupt_line [1])
    );
    X_OR2 \bridge/configuration/interrupt_line<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/interrupt_line[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/interrupt_line[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [4])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<5>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_reg<5> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr [5])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<5>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_latency_tim_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_latency_tim_out[1]/SRNOT )
    );
    X_FF \bridge/configuration/latency_timer_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C283/N39 ),
      .SET (GND),
      .RST (\bridge/conf_latency_tim_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_latency_tim_out [0])
    );
    X_OR2 \bridge/conf_latency_tim_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_latency_tim_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_latency_tim_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/latency_timer_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [9]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C283/N39 ),
      .SET (GND),
      .RST (\bridge/conf_latency_tim_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_latency_tim_out [1])
    );
    X_OR2 \bridge/conf_latency_tim_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_latency_tim_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_latency_tim_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[31]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<30> (
      .I (\bridge/pciu_err_addr_out[30] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [30])
    );
    X_OR2 \bridge/configuration/pci_err_addr<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<31> (
      .I (\bridge/pciu_err_addr_out[31] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [31])
    );
    X_OR2 \bridge/configuration/pci_err_addr<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[23]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<22> (
      .I (\bridge/pciu_err_addr_out[22] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [22])
    );
    X_OR2 \bridge/configuration/pci_err_addr<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<23> (
      .I (\bridge/pciu_err_addr_out[23] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [23])
    );
    X_OR2 \bridge/configuration/pci_err_addr<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<14> (
      .I (\bridge/pciu_err_addr_out[14] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [14])
    );
    X_OR2 \bridge/configuration/pci_err_addr<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<15> (
      .I (\bridge/pciu_err_addr_out[15] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [15])
    );
    X_OR2 \bridge/configuration/pci_err_addr<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/interrupt_line<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/interrupt_line[3]/SRNOT )
    );
    X_FF \bridge/configuration/interrupt_line_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C288/N39 ),
      .SET (GND),
      .RST (\bridge/configuration/interrupt_line[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/interrupt_line [2])
    );
    X_OR2 \bridge/configuration/interrupt_line<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/interrupt_line[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/interrupt_line[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/interrupt_line_reg<3> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C288/N39 ),
      .SET (GND),
      .RST (\bridge/configuration/interrupt_line[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/interrupt_line [3])
    );
    X_OR2 \bridge/configuration/interrupt_line<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/interrupt_line[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/interrupt_line[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_latency_tim_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_latency_tim_out[3]/SRNOT )
    );
    X_FF \bridge/configuration/latency_timer_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [10]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C283/N39 ),
      .SET (GND),
      .RST (\bridge/conf_latency_tim_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_latency_tim_out [2])
    );
    X_OR2 \bridge/conf_latency_tim_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_latency_tim_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_latency_tim_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/latency_timer_reg<3> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [11]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C283/N39 ),
      .SET (GND),
      .RST (\bridge/conf_latency_tim_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_latency_tim_out [3])
    );
    X_OR2 \bridge/conf_latency_tim_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_latency_tim_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_latency_tim_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[25]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<24> (
      .I (\bridge/pciu_err_addr_out[24] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [24])
    );
    X_OR2 \bridge/configuration/pci_err_addr<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<25> (
      .I (\bridge/pciu_err_addr_out[25] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [25])
    );
    X_OR2 \bridge/configuration/pci_err_addr<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<16> (
      .I (\bridge/pciu_err_addr_out[16] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [16])
    );
    X_OR2 \bridge/configuration/pci_err_addr<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<17> (
      .I (\bridge/pciu_err_addr_out[17] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [17])
    );
    X_OR2 \bridge/configuration/pci_err_addr<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/interrupt_line<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/interrupt_line[5]/SRNOT )
    );
    X_FF \bridge/configuration/interrupt_line_reg<4> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C288/N39 ),
      .SET (GND),
      .RST (\bridge/configuration/interrupt_line[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/interrupt_line [4])
    );
    X_OR2 \bridge/configuration/interrupt_line<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/interrupt_line[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/interrupt_line[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/interrupt_line_reg<5> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C288/N39 ),
      .SET (GND),
      .RST (\bridge/configuration/interrupt_line[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/interrupt_line [5])
    );
    X_OR2 \bridge/configuration/interrupt_line<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/interrupt_line[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/interrupt_line[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_latency_tim_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_latency_tim_out[5]/SRNOT )
    );
    X_FF \bridge/configuration/latency_timer_reg<4> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C283/N39 ),
      .SET (GND),
      .RST (\bridge/conf_latency_tim_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_latency_tim_out [4])
    );
    X_OR2 \bridge/conf_latency_tim_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_latency_tim_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_latency_tim_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/latency_timer_reg<5> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C283/N39 ),
      .SET (GND),
      .RST (\bridge/conf_latency_tim_out[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_latency_tim_out [5])
    );
    X_OR2 \bridge/conf_latency_tim_out<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_latency_tim_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_latency_tim_out[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[27]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<26> (
      .I (\bridge/pciu_err_addr_out[26] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [26])
    );
    X_OR2 \bridge/configuration/pci_err_addr<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<27> (
      .I (\bridge/pciu_err_addr_out[27] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [27])
    );
    X_OR2 \bridge/configuration/pci_err_addr<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<18> (
      .I (\bridge/pciu_err_addr_out[18] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [18])
    );
    X_OR2 \bridge/configuration/pci_err_addr<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<19> (
      .I (\bridge/pciu_err_addr_out[19] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [19])
    );
    X_OR2 \bridge/configuration/pci_err_addr<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/SRNOT )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<0>/BYMUX (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [0]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/BYNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[0]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/interrupt_line<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/interrupt_line[7]/SRNOT )
    );
    X_FF \bridge/configuration/interrupt_line_reg<6> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C288/N39 ),
      .SET (GND),
      .RST (\bridge/configuration/interrupt_line[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/interrupt_line [6])
    );
    X_OR2 \bridge/configuration/interrupt_line<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/interrupt_line[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/interrupt_line[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/interrupt_line_reg<7> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C288/N39 ),
      .SET (GND),
      .RST (\bridge/configuration/interrupt_line[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/interrupt_line [7])
    );
    X_OR2 \bridge/configuration/interrupt_line<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/interrupt_line[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/interrupt_line[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/int_prop_en/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/int_prop_en/SRNOT )
    );
    X_FF \bridge/configuration/icr_bit3_0_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C302/N19 ),
      .SET (GND),
      .RST (\bridge/configuration/int_prop_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/int_prop_en )
    );
    X_OR2 \bridge/configuration/int_prop_en/FFY/ASYNC_FF_GSR_OR_137 (
      .I0 (\bridge/configuration/int_prop_en/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/int_prop_en/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_latency_tim_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_latency_tim_out[7]/SRNOT )
    );
    X_FF \bridge/configuration/latency_timer_reg<6> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C283/N39 ),
      .SET (GND),
      .RST (\bridge/conf_latency_tim_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_latency_tim_out [6])
    );
    X_OR2 \bridge/conf_latency_tim_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_latency_tim_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_latency_tim_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/latency_timer_reg<7> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C283/N39 ),
      .SET (GND),
      .RST (\bridge/conf_latency_tim_out[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_latency_tim_out [7])
    );
    X_OR2 \bridge/conf_latency_tim_out<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_latency_tim_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_latency_tim_out[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/error_int_en/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/error_int_en/SRNOT )
    );
    X_FF \bridge/configuration/icr_bit3_0_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C302/N19 ),
      .SET (GND),
      .RST (\bridge/configuration/error_int_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/error_int_en )
    );
    X_OR2 \bridge/configuration/error_int_en/FFY/ASYNC_FF_GSR_OR_138 (
      .I0 (\bridge/configuration/error_int_en/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/error_int_en/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[29]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<28> (
      .I (\bridge/pciu_err_addr_out[28] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [28])
    );
    X_OR2 \bridge/configuration/pci_err_addr<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<29> (
      .I (\bridge/pciu_err_addr_out[29] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [29])
    );
    X_OR2 \bridge/configuration/pci_err_addr<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/perr_int_en/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/perr_int_en/SRNOT )
    );
    X_FF \bridge/configuration/icr_bit3_0_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C302/N19 ),
      .SET (GND),
      .RST (\bridge/configuration/perr_int_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/perr_int_en )
    );
    X_OR2 \bridge/configuration/perr_int_en/FFY/ASYNC_FF_GSR_OR_139 (
      .I0 (\bridge/configuration/perr_int_en/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/perr_int_en/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr1<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr1[21]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [20])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [21])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr1<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr1[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [12])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [13])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/serr_int_en/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/serr_int_en/SRNOT )
    );
    X_FF \bridge/configuration/icr_bit3_0_reg<3> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C302/N19 ),
      .SET (GND),
      .RST (\bridge/configuration/serr_int_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/serr_int_en )
    );
    X_OR2 \bridge/configuration/serr_int_en/FFY/ASYNC_FF_GSR_OR_140 (
      .I0 (\bridge/configuration/serr_int_en/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/serr_int_en/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_ba1_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_ba1_out[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<30> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N19 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba1_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba1_out [18])
    );
    X_OR2 \bridge/conf_pci_ba1_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba1_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba1_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<31> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N19 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba1_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba1_out [19])
    );
    X_OR2 \bridge/conf_pci_ba1_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba1_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba1_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr1<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr1[23]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [22])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [23])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr1<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr1[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [14])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [15])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_ba1_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_ba1_out[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<24> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N19 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba1_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba1_out [12])
    );
    X_OR2 \bridge/conf_pci_ba1_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba1_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba1_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<25> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N19 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba1_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba1_out [13])
    );
    X_OR2 \bridge/conf_pci_ba1_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba1_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba1_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr1<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr1[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [16])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [17])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[1]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<0> (
      .I (\bridge/out_bckp_ad_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [0])
    );
    X_OR2 \bridge/configuration/wb_err_data<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<1> (
      .I (\bridge/out_bckp_ad_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [1])
    );
    X_OR2 \bridge/configuration/wb_err_data<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C120 .INIT = 16'hF0FA;
    X_LUT4 \bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/C120 (
      .ADR0 (\bridge/pci_target_unit/pcit_if_pcir_fifo_data_err_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pcit_if_disconect_wo_data_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy/GROM )
    );
    defparam C19134.INIT = 16'h5000;
    X_LUT4 C19134(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/N64 ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_pcir_fifo_data_err_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy/GROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/pci_target_clock_en/syn129 )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/devs_w_frm_irdy )
    );
    X_INV \bridge/conf_pci_ba1_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_ba1_out[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<26> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N19 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba1_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba1_out [14])
    );
    X_OR2 \bridge/conf_pci_ba1_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba1_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba1_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<27> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N19 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba1_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba1_out [15])
    );
    X_OR2 \bridge/conf_pci_ba1_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba1_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba1_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr1<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr1[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [18])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N54 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr1[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr1 [19])
    );
    X_OR2 \bridge/configuration/pci_base_addr1<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr1[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr1[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[3]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<2> (
      .I (\bridge/out_bckp_ad_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [2])
    );
    X_OR2 \bridge/configuration/wb_err_data<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<3> (
      .I (\bridge/out_bckp_ad_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [3])
    );
    X_OR2 \bridge/configuration/wb_err_data<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/conf_pci_ba1_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_ba1_out[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<28> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N19 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba1_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba1_out [16])
    );
    X_OR2 \bridge/conf_pci_ba1_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba1_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba1_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba1_bit31_12_reg<29> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C286/N19 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba1_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba1_out [17])
    );
    X_OR2 \bridge/conf_pci_ba1_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba1_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba1_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/wb_err_data<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[5]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<4> (
      .I (\bridge/out_bckp_ad_out [4]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [4])
    );
    X_OR2 \bridge/configuration/wb_err_data<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<5> (
      .I (\bridge/out_bckp_ad_out [5]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [5])
    );
    X_OR2 \bridge/configuration/wb_err_data<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [2])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [3])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/wb_err_data<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[7]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<6> (
      .I (\bridge/out_bckp_ad_out [6]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [6])
    );
    X_OR2 \bridge/configuration/wb_err_data<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<7> (
      .I (\bridge/out_bckp_ad_out [7]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [7])
    );
    X_OR2 \bridge/configuration/wb_err_data<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18020.INIT = 16'hCDCC;
    X_LUT4 C18020(
      .ADR0 (syn18863),
      .ADR1 (N12594),
      .ADR2 (N_TRDY),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .O (\syn22225/GROM )
    );
    defparam C18069.INIT = 16'h0004;
    X_LUT4 C18069(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_last_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/posted_write_req ),
      .ADR2 (syn18863),
      .ADR3 (N_TRDY),
      .O (\syn22225/FROM )
    );
    X_BUF \syn22225/YUSED (
      .I (\syn22225/GROM ),
      .O (N12436)
    );
    X_BUF \syn22225/XUSED (
      .I (\syn22225/FROM ),
      .O (syn22225)
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[4]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/wb_err_data<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_err_data[9]/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_data_reg<8> (
      .I (\bridge/out_bckp_ad_out [8]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [8])
    );
    X_OR2 \bridge/configuration/wb_err_data<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/wb_err_data_reg<9> (
      .I (\bridge/out_bckp_ad_out [9]),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/configuration/wb_err_data[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_err_data [9])
    );
    X_OR2 \bridge/configuration/wb_err_data<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/wb_err_data[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_err_data[9]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18200.INIT = 16'h7DBE;
    X_LUT4 C18200(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/inGreyCount [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/inGreyCount [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/outGreyCount [3]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/outGreyCount [2]),
      .O (\syn181402/GROM )
    );
    X_BUF \syn181402/YUSED (
      .I (\syn181402/GROM ),
      .O (syn181402)
    );
    defparam C18112.INIT = 16'hA0A0;
    X_LUT4 C18112(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/GROM )
    );
    defparam C18113.INIT = 16'h33FF;
    X_LUT4 C18113(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_clr ),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg ),
      .O (N12592)
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/GROM ),
      .O (N12378)
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg_reg (
      .I (N12592),
      .CLK (CLK_BUFGPed),
      .CE (N12378),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/FFX/ASYNC_FF_GSR_OR_141 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_rty_exp_reg/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18130.INIT = 16'hDCFF;
    X_LUT4 C18130(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 ),
      .ADR1 (syn18863),
      .ADR2 (syn19064),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/del_write_req ),
      .O (\bridge/wbu_mabort_rec_out/GROM )
    );
    defparam C18134.INIT = 16'h4444;
    X_LUT4 C18134(
      .ADR0 (syn18863),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/S_60/cell0 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wbu_mabort_rec_out/FROM )
    );
    X_INV \bridge/wbu_mabort_rec_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wbu_mabort_rec_out/SRNOT )
    );
    X_BUF \bridge/wbu_mabort_rec_out/YUSED (
      .I (\bridge/wbu_mabort_rec_out/GROM ),
      .O (syn22095)
    );
    X_BUF \bridge/wbu_mabort_rec_out/XUSED (
      .I (\bridge/wbu_mabort_rec_out/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/tabort_ff_in )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/tabort_received_out_reg (
      .I (\bridge/wbu_mabort_rec_out/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/wbu_mabort_rec_out/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wbu_mabort_rec_out )
    );
    X_OR2 \bridge/wbu_mabort_rec_out/FFX/ASYNC_FF_GSR_OR_142 (
      .I0 (\bridge/wbu_mabort_rec_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wbu_mabort_rec_out/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18114.INIT = 16'hBBFF;
    X_LUT4 C18114(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [16]),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/req_comp_pending_sample ),
      .ADR2 (VCC),
      .ADR3 (syn22126),
      .O (\N12380/GROM )
    );
    defparam C18118.INIT = 16'hBBFF;
    X_LUT4 C18118(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [16]),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/req_done_reg ),
      .ADR2 (VCC),
      .ADR3 (syn22126),
      .O (\N12380/FROM )
    );
    X_BUF \N12380/YUSED (
      .I (\N12380/GROM ),
      .O (N12379)
    );
    X_BUF \N12380/XUSED (
      .I (\N12380/FROM ),
      .O (N12380)
    );
    defparam C18203.INIT = 16'h0011;
    X_LUT4 C18203(
      .ADR0 (N12360),
      .ADR1 (syn177324),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_full_out ),
      .O (\N12607/GROM )
    );
    defparam C19449.INIT = 16'hFFFA;
    X_LUT4 C19449(
      .ADR0 (N12360),
      .ADR1 (VCC),
      .ADR2 (syn177324),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_full_out ),
      .O (\N12607/FROM )
    );
    X_BUF \N12607/YUSED (
      .I (\N12607/GROM ),
      .O (\bridge/wishbone_slave_unit/fifos/in_count_en )
    );
    X_BUF \N12607/XUSED (
      .I (\N12607/FROM ),
      .O (N12607)
    );
    defparam C18212.INIT = 16'h505F;
    X_LUT4 C18212(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .O (\syn18930/GROM )
    );
    defparam C19457.INIT = 16'h3030;
    X_LUT4 C19457(
      .ADR0 (VCC),
      .ADR1 (\bridge/out_bckp_frame_out ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (VCC),
      .O (\syn18930/FROM )
    );
    X_BUF \syn18930/YUSED (
      .I (\syn18930/GROM ),
      .O (N12351)
    );
    X_BUF \syn18930/XUSED (
      .I (\syn18930/FROM ),
      .O (syn18930)
    );
    defparam C18116.INIT = 16'h22F2;
    X_LUT4 C18116(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main ),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync_comp_req_pending_out ),
      .ADR3 (syn22096),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/GROM )
    );
    defparam C18117.INIT = 16'hCFCF;
    X_LUT4 C18117(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_clr ),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/comp_done_reg_main ),
      .ADR3 (VCC),
      .O (N12593)
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/GROM ),
      .O (N12381)
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_comp_pending_reg (
      .I (N12593),
      .CLK (CLK_BUFGPed),
      .CE (N12381),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/FFX/ASYNC_FF_GSR_OR_143 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[4]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/raddr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pciw_rallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [4])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[4]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next[4]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C18310.INIT = 16'hEAC0;
    X_LUT4 C18310(
      .ADR0 (syn16919),
      .ADR1 (syn16931),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [29]),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [29]),
      .O (\syn181005/GROM )
    );
    defparam C18368.INIT = 16'hF888;
    X_LUT4 C18368(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [26]),
      .ADR1 (syn16919),
      .ADR2 (syn16931),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [26]),
      .O (\syn181005/FROM )
    );
    X_BUF \syn181005/YUSED (
      .I (\syn181005/GROM ),
      .O (syn120398)
    );
    X_BUF \syn181005/XUSED (
      .I (\syn181005/FROM ),
      .O (syn181005)
    );
    defparam C18070.INIT = 16'h0307;
    X_LUT4 C18070(
      .ADR0 (N_TRDY),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_rdy_out ),
      .ADR2 (N12594),
      .ADR3 (syn18863),
      .O (\N12466/GROM )
    );
    defparam C18090.INIT = 16'h1F0F;
    X_LUT4 C18090(
      .ADR0 (syn18863),
      .ADR1 (N_TRDY),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_burst_out ),
      .O (\N12466/FROM )
    );
    X_BUF \N12466/YUSED (
      .I (\N12466/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/last_load )
    );
    X_BUF \N12466/XUSED (
      .I (\N12466/FROM ),
      .O (N12466)
    );
    defparam C18303.INIT = 16'hF888;
    X_LUT4 C18303(
      .ADR0 (\bridge/configuration/wb_err_addr [30]),
      .ADR1 (\bridge/configuration/C1937 ),
      .ADR2 (\bridge/configuration/wb_err_cs_bit31_24 [30]),
      .ADR3 (\bridge/configuration/C1941 ),
      .O (\syn181040/GROM )
    );
    defparam C18359.INIT = 16'hECA0;
    X_LUT4 C18359(
      .ADR0 (\bridge/configuration/wb_err_addr [27]),
      .ADR1 (\bridge/configuration/C1941 ),
      .ADR2 (\bridge/configuration/C1937 ),
      .ADR3 (\bridge/configuration/wb_err_cs_bit31_24 [27]),
      .O (\syn181040/FROM )
    );
    X_BUF \syn181040/YUSED (
      .I (\syn181040/GROM ),
      .O (syn181196)
    );
    X_BUF \syn181040/XUSED (
      .I (\syn181040/FROM ),
      .O (syn181040)
    );
    defparam C18223.INIT = 16'hFF40;
    X_LUT4 C18223(
      .ADR0 (\bridge/out_bckp_frame_out ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_time_out ),
      .ADR2 (N_GNT),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout ),
      .O (\syn178588/GROM )
    );
    defparam C19460.INIT = 16'hFEFE;
    X_LUT4 C19460(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/timeout ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_last_out ),
      .ADR3 (VCC),
      .O (\syn178588/FROM )
    );
    X_BUF \syn178588/YUSED (
      .I (\syn178588/GROM ),
      .O (syn21738)
    );
    X_BUF \syn178588/XUSED (
      .I (\syn178588/FROM ),
      .O (syn178588)
    );
    defparam C19200.INIT = 16'hCFC0;
    X_LUT4 C19200(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [14]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[14]/GROM )
    );
    defparam C19343.INIT = 16'hFFCC;
    X_LUT4 C19343(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[14]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<14>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[14]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [14])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<14>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[14]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [14])
    );
    defparam C18320.INIT = 16'hEAC0;
    X_LUT4 C18320(
      .ADR0 (\bridge/configuration/C1989 ),
      .ADR1 (\bridge/configuration/C2003 ),
      .ADR2 (\bridge/conf_pci_ba0_out [17]),
      .ADR3 (\bridge/conf_pci_am1_out [17]),
      .O (\syn181092/GROM )
    );
    defparam C18338.INIT = 16'hECA0;
    X_LUT4 C18338(
      .ADR0 (\bridge/configuration/C1989 ),
      .ADR1 (\bridge/configuration/C2003 ),
      .ADR2 (\bridge/conf_pci_am1_out [16]),
      .ADR3 (\bridge/conf_pci_ba0_out [16]),
      .O (\syn181092/FROM )
    );
    X_BUF \syn181092/YUSED (
      .I (\syn181092/GROM ),
      .O (syn181143)
    );
    X_BUF \syn181092/XUSED (
      .I (\syn181092/FROM ),
      .O (syn181092)
    );
    defparam C18304.INIT = 16'hEAC0;
    X_LUT4 C18304(
      .ADR0 (\bridge/configuration/C2003 ),
      .ADR1 (\bridge/configuration/C1935 ),
      .ADR2 (\bridge/configuration/wb_err_data [30]),
      .ADR3 (\bridge/conf_pci_ba0_out [18]),
      .O (\syn181039/GROM )
    );
    defparam C18360.INIT = 16'hECA0;
    X_LUT4 C18360(
      .ADR0 (\bridge/configuration/C2003 ),
      .ADR1 (\bridge/configuration/wb_err_data [27]),
      .ADR2 (\bridge/conf_pci_ba0_out [15]),
      .ADR3 (\bridge/configuration/C1935 ),
      .O (\syn181039/FROM )
    );
    X_BUF \syn181039/YUSED (
      .I (\syn181039/GROM ),
      .O (syn181195)
    );
    X_BUF \syn181039/XUSED (
      .I (\syn181039/FROM ),
      .O (syn181039)
    );
    defparam C19201.INIT = 16'hFC0C;
    X_LUT4 C19201(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_addr_out [15]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[0]/GROM )
    );
    defparam C19212.INIT = 16'hFC0C;
    X_LUT4 C19212(
      .ADR0 (VCC),
      .ADR1 (\bridge/in_reg_cbe_out [0]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_bc_out [0]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[0]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out<0>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[0]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [15])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out<0>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[0]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out [0])
    );
    defparam C19041.INIT = 16'h0003;
    X_LUT4 C19041(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_wbm_if/vmaddr_r [1]),
      .ADR2 (\CRT/ssvga_wbm_if/vmaddr_r [0]),
      .ADR3 (\CRT/ssvga_wbm_if/vmaddr_r [16]),
      .O (\CRT/ssvga_wbm_if/N1531/GROM )
    );
    defparam C19110.INIT = 16'h00FF;
    X_LUT4 C19110(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/vmaddr_r [16]),
      .O (N12635)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C19/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C18/C1/O ),
      .I1 (N12635),
      .O (\CRT/ssvga_wbm_if/N1531/XORF )
    );
    X_BUF \CRT/ssvga_wbm_if/N1531/YUSED (
      .I (\CRT/ssvga_wbm_if/N1531/GROM ),
      .O (syn179376)
    );
    X_BUF \CRT/ssvga_wbm_if/N1531/XUSED (
      .I (\CRT/ssvga_wbm_if/N1531/XORF ),
      .O (\CRT/ssvga_wbm_if/N1531 )
    );
    defparam C18225.INIT = 16'h0001;
    X_LUT4 C18225(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [3]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [2]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [4]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [5]),
      .O (\syn181347/GROM )
    );
    X_BUF \syn181347/YUSED (
      .I (\syn181347/GROM ),
      .O (syn181347)
    );
    defparam C18161.INIT = 16'hC03F;
    X_LUT4 C18161(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [19]),
      .ADR2 (syn24500),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [19]),
      .O (\syn17084/GROM )
    );
    defparam C19569.INIT = 16'hC000;
    X_LUT4 C19569(
      .ADR0 (VCC),
      .ADR1 (syn24500),
      .ADR2 (syn177629),
      .ADR3 (syn16936),
      .O (\syn17084/FROM )
    );
    X_BUF \syn17084/YUSED (
      .I (\syn17084/GROM ),
      .O (syn176967)
    );
    X_BUF \syn17084/XUSED (
      .I (\syn17084/FROM ),
      .O (syn17084)
    );
    defparam C19202.INIT = 16'h0008;
    X_LUT4 C19202(
      .ADR0 (syn19713),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .ADR2 (\bridge/pci_target_unit/del_sync_bc_out [0]),
      .ADR3 (syn19710),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[0]/GROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out<0>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out[0]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out [0])
    );
    defparam C19042.INIT = 16'h0001;
    X_LUT4 C19042(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [6]),
      .ADR1 (\CRT/ssvga_wbm_if/vmaddr_r [7]),
      .ADR2 (\CRT/ssvga_wbm_if/vmaddr_r [8]),
      .ADR3 (\CRT/ssvga_wbm_if/vmaddr_r [9]),
      .O (\syn179378/GROM )
    );
    X_BUF \syn179378/YUSED (
      .I (\syn179378/GROM ),
      .O (syn179378)
    );
    defparam C18402.INIT = 16'hEAC0;
    X_LUT4 C18402(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_data_out [24]),
      .ADR2 (syn20493),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [24]),
      .O (\syn180806/GROM )
    );
    defparam C18434.INIT = 16'hF888;
    X_LUT4 C18434(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [22]),
      .ADR2 (syn20493),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [22]),
      .O (\syn180806/FROM )
    );
    X_BUF \syn180806/YUSED (
      .I (\syn180806/GROM ),
      .O (syn180899)
    );
    X_BUF \syn180806/XUSED (
      .I (\syn180806/FROM ),
      .O (syn180806)
    );
    defparam C18314.INIT = 16'hECA0;
    X_LUT4 C18314(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [29]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_data_out [29]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (syn20493),
      .O (\syn181107/GROM )
    );
    defparam C18332.INIT = 16'hECA0;
    X_LUT4 C18332(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [28]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_data_out [28]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .O (\syn181107/FROM )
    );
    X_BUF \syn181107/YUSED (
      .I (\syn181107/GROM ),
      .O (syn181158)
    );
    X_BUF \syn181107/XUSED (
      .I (\syn181107/FROM ),
      .O (syn181107)
    );
    defparam C19211.INIT = 16'hF8FF;
    X_LUT4 C19211(
      .ADR0 (\bridge/pci_target_unit/del_sync_bc_out [2]),
      .ADR1 (\bridge/pci_target_unit/del_sync_burst_out ),
      .ADR2 (\bridge/pci_target_unit/del_sync_bc_out [3]),
      .ADR3 (\bridge/pci_target_unit/del_sync_bc_out [1]),
      .O (\syn19708/GROM )
    );
    X_BUF \syn19708/YUSED (
      .I (\syn19708/GROM ),
      .O (syn19708)
    );
    defparam C19203.INIT = 16'h5050;
    X_LUT4 C19203(
      .ADR0 (ERR_I),
      .ADR1 (VCC),
      .ADR2 (ACK_I),
      .ADR3 (VCC),
      .O (\syn19562/GROM )
    );
    defparam C19254.INIT = 16'h5A5A;
    X_LUT4 C19254(
      .ADR0 (ACK_I),
      .ADR1 (VCC),
      .ADR2 (ERR_I),
      .ADR3 (VCC),
      .O (\syn19562/FROM )
    );
    X_BUF \syn19562/YUSED (
      .I (\syn19562/GROM ),
      .O (syn19713)
    );
    X_BUF \syn19562/XUSED (
      .I (\syn19562/FROM ),
      .O (syn19562)
    );
    defparam C19043.INIT = 16'h0001;
    X_LUT4 C19043(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [3]),
      .ADR1 (\CRT/ssvga_wbm_if/vmaddr_r [5]),
      .ADR2 (\CRT/ssvga_wbm_if/vmaddr_r [2]),
      .ADR3 (\CRT/ssvga_wbm_if/vmaddr_r [4]),
      .O (\syn179377/GROM )
    );
    X_BUF \syn179377/YUSED (
      .I (\syn179377/GROM ),
      .O (syn179377)
    );
    defparam C18411.INIT = 16'hEC00;
    X_LUT4 C18411(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/configuration/C1953 ),
      .ADR2 (\bridge/conf_wb_ba1_out [12]),
      .ADR3 (\bridge/conf_wb_am1_out [12]),
      .O (\syn60043/GROM )
    );
    defparam C19968.INIT = 16'hA5FF;
    X_LUT4 C19968(
      .ADR0 (\bridge/conf_wb_ba1_out [12]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [24]),
      .ADR3 (\bridge/conf_wb_am1_out [12]),
      .O (\syn60043/FROM )
    );
    X_BUF \syn60043/YUSED (
      .I (\syn60043/GROM ),
      .O (syn21325)
    );
    X_BUF \syn60043/XUSED (
      .I (\syn60043/FROM ),
      .O (syn60043)
    );
    defparam C18323.INIT = 16'hC8C0;
    X_LUT4 C18323(
      .ADR0 (\bridge/conf_wb_ba1_out [17]),
      .ADR1 (\bridge/conf_wb_am1_out [17]),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/configuration/C1955 ),
      .O (\syn60048/GROM )
    );
    defparam C19971.INIT = 16'hF55F;
    X_LUT4 C19971(
      .ADR0 (\bridge/conf_wb_am1_out [17]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [29]),
      .ADR3 (\bridge/conf_wb_ba1_out [17]),
      .O (\syn60048/FROM )
    );
    X_BUF \syn60048/YUSED (
      .I (\syn60048/GROM ),
      .O (syn21531)
    );
    X_BUF \syn60048/XUSED (
      .I (\syn60048/FROM ),
      .O (syn60048)
    );
    defparam C18147.INIT = 16'h6006;
    X_LUT4 C18147(
      .ADR0 (\bridge/wishbone_slave_unit/del_sync_addr_out [7]),
      .ADR1 (syn60030),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync_addr_out [8]),
      .O (\syn17119/GROM )
    );
    defparam C19577.INIT = 16'h4000;
    X_LUT4 C19577(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR1 (syn60030),
      .ADR2 (syn17772),
      .ADR3 (syn59978),
      .O (\syn17119/FROM )
    );
    X_BUF \syn17119/YUSED (
      .I (\syn17119/GROM ),
      .O (syn181509)
    );
    X_BUF \syn17119/XUSED (
      .I (\syn17119/FROM ),
      .O (syn17119)
    );
    defparam C19060.INIT = 16'h0A0A;
    X_LUT4 C19060(
      .ADR0 (\CRT/pal_pix_dat [11]),
      .ADR1 (VCC),
      .ADR2 (\CRT/drive_blank_reg ),
      .ADR3 (VCC),
      .O (\rgb_int[10]/GROM )
    );
    defparam C19061.INIT = 16'h5050;
    X_LUT4 C19061(
      .ADR0 (\CRT/drive_blank_reg ),
      .ADR1 (VCC),
      .ADR2 (\CRT/pal_pix_dat [10]),
      .ADR3 (VCC),
      .O (\rgb_int[10]/FROM )
    );
    X_BUF \rgb_int<10>/YUSED (
      .I (\rgb_int[10]/GROM ),
      .O (rgb_int[11])
    );
    X_BUF \rgb_int<10>/XUSED (
      .I (\rgb_int[10]/FROM ),
      .O (rgb_int[10])
    );
    defparam C18180.INIT = 16'h1000;
    X_LUT4 C18180(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [0]),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .ADR2 (\CRT/ssvga_wbm_if/S_41/cell0 ),
      .ADR3 (syn177324),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C707/GROM )
    );
    defparam C19979.INIT = 16'h00A0;
    X_LUT4 C19979(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [0]),
      .ADR3 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [1]),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C707/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/C707/YUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/C707/GROM ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/C707/XUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/C707/FROM ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/C707 )
    );
    defparam C19213.INIT = 16'hF0CC;
    X_LUT4 C19213(
      .ADR0 (VCC),
      .ADR1 (\bridge/in_reg_cbe_out [1]),
      .ADR2 (\bridge/pci_target_unit/pcit_if_bc_out [1]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[2]/GROM )
    );
    defparam C19214.INIT = 16'hFC0C;
    X_LUT4 C19214(
      .ADR0 (VCC),
      .ADR1 (\bridge/in_reg_cbe_out [2]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_bc_out [2]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[2]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out<2>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[2]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out [1])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out<2>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[2]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out [2])
    );
    defparam C18501.INIT = 16'hEAC0;
    X_LUT4 C18501(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (\bridge/configuration/wb_err_addr [18]),
      .ADR2 (\bridge/configuration/C1937 ),
      .ADR3 (\bridge/configuration/wb_err_data [18]),
      .O (\syn180469/GROM )
    );
    defparam C18548.INIT = 16'hF888;
    X_LUT4 C18548(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (\bridge/configuration/wb_err_data [15]),
      .ADR2 (\bridge/configuration/C1937 ),
      .ADR3 (\bridge/configuration/wb_err_addr [15]),
      .O (\syn180469/FROM )
    );
    X_BUF \syn180469/YUSED (
      .I (\syn180469/GROM ),
      .O (syn180610)
    );
    X_BUF \syn180469/XUSED (
      .I (\syn180469/FROM ),
      .O (syn180469)
    );
    defparam C18405.INIT = 16'hF888;
    X_LUT4 C18405(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/configuration/pci_err_addr [24]),
      .ADR2 (\bridge/configuration/C1973 ),
      .ADR3 (\bridge/configuration/pci_err_cs_bit31_24 [24]),
      .O (\syn16983/GROM )
    );
    defparam C18698.INIT = 16'hC0C0;
    X_LUT4 C18698(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/C1971 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (VCC),
      .O (\syn16983/FROM )
    );
    X_BUF \syn16983/YUSED (
      .I (\syn16983/GROM ),
      .O (syn180887)
    );
    X_BUF \syn16983/XUSED (
      .I (\syn16983/FROM ),
      .O (syn16983)
    );
    defparam C18341.INIT = 16'hCC80;
    X_LUT4 C18341(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/conf_wb_am1_out [16]),
      .ADR2 (\bridge/conf_wb_ba1_out [16]),
      .ADR3 (\bridge/configuration/C1953 ),
      .O (\syn60047/GROM )
    );
    defparam C19972.INIT = 16'h99FF;
    X_LUT4 C19972(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [28]),
      .ADR1 (\bridge/conf_wb_ba1_out [16]),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_wb_am1_out [16]),
      .O (\syn60047/FROM )
    );
    X_BUF \syn60047/YUSED (
      .I (\syn60047/GROM ),
      .O (syn21490)
    );
    X_BUF \syn60047/XUSED (
      .I (\syn60047/FROM ),
      .O (syn60047)
    );
    defparam C18085.INIT = 16'hC888;
    X_LUT4 C18085(
      .ADR0 (syn18863),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR2 (syn181624),
      .ADR3 (syn22184),
      .O (\syn181605/GROM )
    );
    defparam C18093.INIT = 16'h0004;
    X_LUT4 C18093(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [3]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/del_read_req ),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [4]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [2]),
      .O (\syn181605/FROM )
    );
    X_BUF \syn181605/YUSED (
      .I (\syn181605/GROM ),
      .O (syn22189)
    );
    X_BUF \syn181605/XUSED (
      .I (\syn181605/FROM ),
      .O (syn181605)
    );
    defparam C19150.INIT = 16'hF000;
    X_LUT4 C19150(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn24519),
      .ADR3 (syn24524),
      .O (\bridge/pci_target_unit/pci_target_sm/ad_en_w/GROM )
    );
    defparam C19153.INIT = 16'hF2F2;
    X_LUT4 C19153(
      .ADR0 (syn17093),
      .ADR1 (\bridge/in_reg_cbe_out [0]),
      .ADR2 (syn24519),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/pci_target_sm/ad_en_w/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/ad_en_w/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/ad_en_w/GROM ),
      .O (syn17035)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/ad_en_w/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/ad_en_w/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/ad_en_w )
    );
    defparam C19070.INIT = 16'h0003;
    X_LUT4 C19070(
      .ADR0 (VCC),
      .ADR1 (syn177321),
      .ADR2 (syn177319),
      .ADR3 (syn177320),
      .O (\CRT/ssvga_fifo/S_43/cell0/GROM )
    );
    X_BUF \CRT/ssvga_fifo/S_43/cell0/YUSED (
      .I (\CRT/ssvga_fifo/S_43/cell0/GROM ),
      .O (\CRT/ssvga_fifo/S_43/cell0 )
    );
    defparam C19062.INIT = 16'h3300;
    X_LUT4 C19062(
      .ADR0 (VCC),
      .ADR1 (\CRT/drive_blank_reg ),
      .ADR2 (VCC),
      .ADR3 (\CRT/pal_pix_dat [9]),
      .O (\rgb_int[8]/GROM )
    );
    defparam C19063.INIT = 16'h3300;
    X_LUT4 C19063(
      .ADR0 (VCC),
      .ADR1 (\CRT/drive_blank_reg ),
      .ADR2 (VCC),
      .ADR3 (\CRT/pal_pix_dat [8]),
      .O (\rgb_int[8]/FROM )
    );
    X_BUF \rgb_int<8>/YUSED (
      .I (\rgb_int[8]/GROM ),
      .O (rgb_int[9])
    );
    X_BUF \rgb_int<8>/XUSED (
      .I (\rgb_int[8]/FROM ),
      .O (rgb_int[8])
    );
    defparam C18422.INIT = 16'hECA0;
    X_LUT4 C18422(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/configuration/pci_err_data [23]),
      .ADR2 (\bridge/configuration/pci_err_addr [23]),
      .ADR3 (\bridge/configuration/C1967 ),
      .O (\syn180794/GROM )
    );
    defparam C18437.INIT = 16'hECA0;
    X_LUT4 C18437(
      .ADR0 (\bridge/configuration/pci_err_data [22]),
      .ADR1 (\bridge/configuration/pci_err_addr [22]),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (\bridge/configuration/C1971 ),
      .O (\syn180794/FROM )
    );
    X_BUF \syn180794/YUSED (
      .I (\syn180794/GROM ),
      .O (syn180844)
    );
    X_BUF \syn180794/XUSED (
      .I (\syn180794/FROM ),
      .O (syn180794)
    );
    defparam C18406.INIT = 16'hF888;
    X_LUT4 C18406(
      .ADR0 (\bridge/configuration/pci_err_data [24]),
      .ADR1 (\bridge/configuration/C1967 ),
      .ADR2 (\bridge/configuration/C1941 ),
      .ADR3 (\bridge/configuration/wb_err_cs_bit31_24 [24]),
      .O (\syn17017/GROM )
    );
    defparam C18858.INIT = 16'hC0C0;
    X_LUT4 C18858(
      .ADR0 (VCC),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1941 ),
      .ADR3 (VCC),
      .O (\syn17017/FROM )
    );
    X_BUF \syn17017/YUSED (
      .I (\syn17017/GROM ),
      .O (syn180886)
    );
    X_BUF \syn17017/XUSED (
      .I (\syn17017/FROM ),
      .O (syn17017)
    );
    defparam C17630.INIT = 16'h9009;
    X_LUT4 C17630(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [1]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [2]),
      .O (\syn182602/GROM )
    );
    defparam C17649.INIT = 16'h7BDE;
    X_LUT4 C17649(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [1]),
      .O (\syn182602/FROM )
    );
    X_BUF \syn182602/YUSED (
      .I (\syn182602/GROM ),
      .O (syn182642)
    );
    X_BUF \syn182602/XUSED (
      .I (\syn182602/FROM ),
      .O (syn182602)
    );
    defparam C18503.INIT = 16'hF888;
    X_LUT4 C18503(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [18]),
      .ADR1 (\bridge/configuration/C1987 ),
      .ADR2 (\bridge/configuration/C1989 ),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [18]),
      .O (\syn180467/GROM )
    );
    defparam C18550.INIT = 16'hECA0;
    X_LUT4 C18550(
      .ADR0 (\bridge/configuration/C1989 ),
      .ADR1 (\bridge/configuration/C1987 ),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [15]),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [15]),
      .O (\syn180467/FROM )
    );
    X_BUF \syn180467/YUSED (
      .I (\syn180467/GROM ),
      .O (syn180608)
    );
    X_BUF \syn180467/XUSED (
      .I (\syn180467/FROM ),
      .O (syn180467)
    );
    defparam C18407.INIT = 16'hEAC0;
    X_LUT4 C18407(
      .ADR0 (\bridge/configuration/wb_err_addr [24]),
      .ADR1 (\bridge/configuration/wb_err_data [24]),
      .ADR2 (\bridge/configuration/C1935 ),
      .ADR3 (\bridge/configuration/C1937 ),
      .O (\syn180843/GROM )
    );
    defparam C18423.INIT = 16'hF888;
    X_LUT4 C18423(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (\bridge/configuration/wb_err_data [23]),
      .ADR2 (\bridge/configuration/C1937 ),
      .ADR3 (\bridge/configuration/wb_err_addr [23]),
      .O (\syn180843/FROM )
    );
    X_BUF \syn180843/YUSED (
      .I (\syn180843/GROM ),
      .O (syn180885)
    );
    X_BUF \syn180843/XUSED (
      .I (\syn180843/FROM ),
      .O (syn180843)
    );
    defparam C18335.INIT = 16'hF888;
    X_LUT4 C18335(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/configuration/pci_err_addr [28]),
      .ADR2 (\bridge/configuration/C1973 ),
      .ADR3 (\bridge/configuration/pci_err_cs_bit31_24 [28]),
      .O (\syn180939/GROM )
    );
    defparam C18388.INIT = 16'hEAC0;
    X_LUT4 C18388(
      .ADR0 (\bridge/configuration/pci_err_addr [25]),
      .ADR1 (\bridge/configuration/pci_err_cs_bit31_24 [25]),
      .ADR2 (\bridge/configuration/C1973 ),
      .ADR3 (\bridge/configuration/C1971 ),
      .O (\syn180939/FROM )
    );
    X_BUF \syn180939/YUSED (
      .I (\syn180939/GROM ),
      .O (syn181095)
    );
    X_BUF \syn180939/XUSED (
      .I (\syn180939/FROM ),
      .O (syn180939)
    );
    defparam C17631.INIT = 16'h9009;
    X_LUT4 C17631(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [4]),
      .O (\syn182601/GROM )
    );
    defparam C17650.INIT = 16'h7DBE;
    X_LUT4 C17650(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_addr [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [3]),
      .O (\syn182601/FROM )
    );
    X_BUF \syn182601/YUSED (
      .I (\syn182601/GROM ),
      .O (syn182641)
    );
    X_BUF \syn182601/XUSED (
      .I (\syn182601/FROM ),
      .O (syn182601)
    );
    defparam C19064.INIT = 16'h5500;
    X_LUT4 C19064(
      .ADR0 (\CRT/drive_blank_reg ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/pal_pix_dat [7]),
      .O (\rgb_int[6]/GROM )
    );
    defparam C19065.INIT = 16'h0C0C;
    X_LUT4 C19065(
      .ADR0 (VCC),
      .ADR1 (\CRT/pal_pix_dat [6]),
      .ADR2 (\CRT/drive_blank_reg ),
      .ADR3 (VCC),
      .O (\rgb_int[6]/FROM )
    );
    X_BUF \rgb_int<6>/YUSED (
      .I (\rgb_int[6]/GROM ),
      .O (rgb_int[7])
    );
    X_BUF \rgb_int<6>/XUSED (
      .I (\rgb_int[6]/FROM ),
      .O (rgb_int[6])
    );
    defparam C19056.INIT = 16'h00CC;
    X_LUT4 C19056(
      .ADR0 (VCC),
      .ADR1 (\CRT/pal_pix_dat [15]),
      .ADR2 (VCC),
      .ADR3 (\CRT/drive_blank_reg ),
      .O (\rgb_int[14]/GROM )
    );
    defparam C19057.INIT = 16'h2222;
    X_LUT4 C19057(
      .ADR0 (\CRT/pal_pix_dat [14]),
      .ADR1 (\CRT/drive_blank_reg ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\rgb_int[14]/FROM )
    );
    X_BUF \rgb_int<14>/YUSED (
      .I (\rgb_int[14]/GROM ),
      .O (rgb_int[15])
    );
    X_BUF \rgb_int<14>/XUSED (
      .I (\rgb_int[14]/FROM ),
      .O (rgb_int[14])
    );
    defparam C18600.INIT = 16'hAA88;
    X_LUT4 C18600(
      .ADR0 (syn181260),
      .ADR1 (syn180322),
      .ADR2 (VCC),
      .ADR3 (syn180321),
      .O (\syn20874/GROM )
    );
    X_BUF \syn20874/YUSED (
      .I (\syn20874/GROM ),
      .O (syn20874)
    );
    defparam C18504.INIT = 16'hECA0;
    X_LUT4 C18504(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [18]),
      .ADR1 (syn17063),
      .ADR2 (\bridge/configuration/C1951 ),
      .ADR3 (syn60110),
      .O (\syn180466/GROM )
    );
    defparam C18551.INIT = 16'hEAC0;
    X_LUT4 C18551(
      .ADR0 (syn60110),
      .ADR1 (\bridge/configuration/C1951 ),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [15]),
      .ADR3 (syn17066),
      .O (\syn180466/FROM )
    );
    X_BUF \syn180466/YUSED (
      .I (\syn180466/GROM ),
      .O (syn180607)
    );
    X_BUF \syn180466/XUSED (
      .I (\syn180466/FROM ),
      .O (syn180466)
    );
    defparam C18440.INIT = 16'hECA0;
    X_LUT4 C18440(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [22]),
      .ADR1 (\bridge/configuration/pci_tran_addr1 [22]),
      .ADR2 (\bridge/configuration/C1989 ),
      .ADR3 (\bridge/configuration/C1987 ),
      .O (\syn180658/GROM )
    );
    defparam C18488.INIT = 16'hEAC0;
    X_LUT4 C18488(
      .ADR0 (\bridge/configuration/C1987 ),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [19]),
      .ADR2 (\bridge/configuration/C1989 ),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [19]),
      .O (\syn180658/FROM )
    );
    X_BUF \syn180658/YUSED (
      .I (\syn180658/GROM ),
      .O (syn180791)
    );
    X_BUF \syn180658/XUSED (
      .I (\syn180658/FROM ),
      .O (syn180658)
    );
    defparam C18432.INIT = 16'hEAC0;
    X_LUT4 C18432(
      .ADR0 (syn136386),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [22]),
      .ADR2 (syn136384),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [22]),
      .O (\syn180763/GROM )
    );
    defparam C18448.INIT = 16'hECA0;
    X_LUT4 C18448(
      .ADR0 (syn136384),
      .ADR1 (\bridge/pci_target_unit/fifos_pcir_data_out [21]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [21]),
      .ADR3 (syn136386),
      .O (\syn180763/FROM )
    );
    X_BUF \syn180763/YUSED (
      .I (\syn180763/GROM ),
      .O (syn180809)
    );
    X_BUF \syn180763/XUSED (
      .I (\syn180763/FROM ),
      .O (syn180763)
    );
    defparam C18424.INIT = 16'hEAC0;
    X_LUT4 C18424(
      .ADR0 (\bridge/configuration/C2003 ),
      .ADR1 (\bridge/configuration/config_addr[23] ),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/configuration/pci_base_addr0 [23]),
      .O (\syn180792/GROM )
    );
    defparam C18439.INIT = 16'hEAC0;
    X_LUT4 C18439(
      .ADR0 (\bridge/configuration/C1929 ),
      .ADR1 (\bridge/configuration/pci_base_addr0 [22]),
      .ADR2 (\bridge/configuration/C2003 ),
      .ADR3 (\bridge/configuration/config_addr[22] ),
      .O (\syn180792/FROM )
    );
    X_BUF \syn180792/YUSED (
      .I (\syn180792/GROM ),
      .O (syn180842)
    );
    X_BUF \syn180792/XUSED (
      .I (\syn180792/FROM ),
      .O (syn180792)
    );
    defparam C18336.INIT = 16'hF888;
    X_LUT4 C18336(
      .ADR0 (\bridge/configuration/wb_err_cs_bit31_24 [28]),
      .ADR1 (\bridge/configuration/C1941 ),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (\bridge/configuration/pci_err_data [28]),
      .O (\syn180938/GROM )
    );
    defparam C18389.INIT = 16'hF888;
    X_LUT4 C18389(
      .ADR0 (\bridge/configuration/C1941 ),
      .ADR1 (\bridge/configuration/wb_err_cs_bit31_24 [25]),
      .ADR2 (\bridge/configuration/pci_err_data [25]),
      .ADR3 (\bridge/configuration/C1967 ),
      .O (\syn180938/FROM )
    );
    X_BUF \syn180938/YUSED (
      .I (\syn180938/GROM ),
      .O (syn181094)
    );
    X_BUF \syn180938/XUSED (
      .I (\syn180938/FROM ),
      .O (syn180938)
    );
    defparam C18280.INIT = 16'hF888;
    X_LUT4 C18280(
      .ADR0 (\bridge/configuration/C1941 ),
      .ADR1 (\bridge/configuration/wb_err_cs_bit31_24 [31]),
      .ADR2 (\bridge/configuration/pci_err_data [31]),
      .ADR3 (\bridge/configuration/C1967 ),
      .O (\syn181145/GROM )
    );
    defparam C18318.INIT = 16'hF888;
    X_LUT4 C18318(
      .ADR0 (\bridge/configuration/pci_err_data [29]),
      .ADR1 (\bridge/configuration/C1967 ),
      .ADR2 (\bridge/configuration/C1941 ),
      .ADR3 (\bridge/configuration/wb_err_cs_bit31_24 [29]),
      .O (\syn181145/FROM )
    );
    X_BUF \syn181145/YUSED (
      .I (\syn181145/GROM ),
      .O (syn181251)
    );
    X_BUF \syn181145/XUSED (
      .I (\syn181145/FROM ),
      .O (syn181145)
    );
    defparam C17720.INIT = 16'h9009;
    X_LUT4 C17720(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [4]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [4]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [5]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [5]),
      .O (\syn182473/GROM )
    );
    defparam C17724.INIT = 16'h6FF6;
    X_LUT4 C17724(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [4]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [4]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [5]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [5]),
      .O (\syn182473/FROM )
    );
    X_BUF \syn182473/YUSED (
      .I (\syn182473/GROM ),
      .O (syn182484)
    );
    X_BUF \syn182473/XUSED (
      .I (\syn182473/FROM ),
      .O (syn182473)
    );
    defparam C17640.INIT = 16'h8421;
    X_LUT4 C17640(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [1]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [2]),
      .O (\syn182628/GROM )
    );
    X_BUF \syn182628/YUSED (
      .I (\syn182628/GROM ),
      .O (syn182628)
    );
    defparam C17616.INIT = 16'h8421;
    X_LUT4 C17616(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [1]),
      .O (\syn182663/GROM )
    );
    defparam C17625.INIT = 16'h9009;
    X_LUT4 C17625(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [2]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [1]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [1]),
      .O (\syn182663/FROM )
    );
    X_BUF \syn182663/YUSED (
      .I (\syn182663/GROM ),
      .O (syn182680)
    );
    X_BUF \syn182663/XUSED (
      .I (\syn182663/FROM ),
      .O (syn182663)
    );
    defparam C19137.INIT = 16'hECEC;
    X_LUT4 C19137(
      .ADR0 (syn24524),
      .ADR1 (syn17093),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/N59 ),
      .ADR3 (VCC),
      .O (\syn178884/GROM )
    );
    defparam C19310.INIT = 16'hAA88;
    X_LUT4 C19310(
      .ADR0 (syn178883),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/N59 ),
      .ADR2 (VCC),
      .ADR3 (syn19397),
      .O (\syn178884/FROM )
    );
    X_BUF \syn178884/YUSED (
      .I (\syn178884/GROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/devs_w )
    );
    X_BUF \syn178884/XUSED (
      .I (\syn178884/FROM ),
      .O (syn178884)
    );
    defparam C19073.INIT = 16'hB333;
    X_LUT4 C19073(
      .ADR0 (\bridge/in_reg_cbe_out [1]),
      .ADR1 (\bridge/in_reg_cbe_out [0]),
      .ADR2 (\bridge/in_reg_cbe_out [3]),
      .ADR3 (\bridge/in_reg_cbe_out [2]),
      .O (\bridge/pci_target_unit/pci_target_if/n_1317/GROM )
    );
    defparam C19075.INIT = 16'h80A0;
    X_LUT4 C19075(
      .ADR0 (\bridge/in_reg_cbe_out [0]),
      .ADR1 (\bridge/in_reg_cbe_out [3]),
      .ADR2 (\bridge/in_reg_cbe_out [1]),
      .ADR3 (\bridge/in_reg_cbe_out [2]),
      .O (\bridge/pci_target_unit/pci_target_if/n_1317/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_if/n_1317/YUSED (
      .I (\bridge/pci_target_unit/pci_target_if/n_1317/GROM ),
      .O (\bridge/pci_target_unit/pci_target_if/n_1352 )
    );
    X_BUF \bridge/pci_target_unit/pci_target_if/n_1317/XUSED (
      .I (\bridge/pci_target_unit/pci_target_if/n_1317/FROM ),
      .O (\bridge/pci_target_unit/pci_target_if/n_1317 )
    );
    defparam C18441.INIT = 16'hEAC0;
    X_LUT4 C18441(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (syn17059),
      .ADR2 (syn60110),
      .ADR3 (\bridge/configuration/wb_tran_addr1 [22]),
      .O (\syn180657/GROM )
    );
    defparam C18489.INIT = 16'hF888;
    X_LUT4 C18489(
      .ADR0 (syn60110),
      .ADR1 (syn17062),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [19]),
      .ADR3 (\bridge/configuration/C1951 ),
      .O (\syn180657/FROM )
    );
    X_BUF \syn180657/YUSED (
      .I (\syn180657/GROM ),
      .O (syn180790)
    );
    X_BUF \syn180657/XUSED (
      .I (\syn180657/FROM ),
      .O (syn180657)
    );
    defparam C18337.INIT = 16'hF888;
    X_LUT4 C18337(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (\bridge/configuration/wb_err_data [28]),
      .ADR2 (\bridge/configuration/wb_err_addr [28]),
      .ADR3 (\bridge/configuration/C1937 ),
      .O (\syn180937/GROM )
    );
    defparam C18390.INIT = 16'hF888;
    X_LUT4 C18390(
      .ADR0 (\bridge/configuration/C1937 ),
      .ADR1 (\bridge/configuration/wb_err_addr [25]),
      .ADR2 (\bridge/configuration/C1935 ),
      .ADR3 (\bridge/configuration/wb_err_data [25]),
      .O (\syn180937/FROM )
    );
    X_BUF \syn180937/YUSED (
      .I (\syn180937/GROM ),
      .O (syn181093)
    );
    X_BUF \syn180937/XUSED (
      .I (\syn180937/FROM ),
      .O (syn180937)
    );
    defparam C18281.INIT = 16'hF888;
    X_LUT4 C18281(
      .ADR0 (\bridge/configuration/C1937 ),
      .ADR1 (\bridge/configuration/wb_err_addr [31]),
      .ADR2 (\bridge/configuration/C1935 ),
      .ADR3 (\bridge/configuration/wb_err_data [31]),
      .O (\syn181144/GROM )
    );
    defparam C18319.INIT = 16'hEAC0;
    X_LUT4 C18319(
      .ADR0 (\bridge/configuration/wb_err_data [29]),
      .ADR1 (\bridge/configuration/C1937 ),
      .ADR2 (\bridge/configuration/wb_err_addr [29]),
      .ADR3 (\bridge/configuration/C1935 ),
      .O (\syn181144/FROM )
    );
    X_BUF \syn181144/YUSED (
      .I (\syn181144/GROM ),
      .O (syn181250)
    );
    X_BUF \syn181144/XUSED (
      .I (\syn181144/FROM ),
      .O (syn181144)
    );
    defparam C18273.INIT = 16'hE0C0;
    X_LUT4 C18273(
      .ADR0 (\bridge/conf_pci_ba0_out [19]),
      .ADR1 (syn120402),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn16929),
      .O (\syn20872/GROM )
    );
    defparam C18594.INIT = 16'h8080;
    X_LUT4 C18594(
      .ADR0 (syn16929),
      .ADR1 (\bridge/configuration/pci_base_addr0 [12]),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (VCC),
      .O (\syn20872/FROM )
    );
    X_BUF \syn20872/YUSED (
      .I (\syn20872/GROM ),
      .O (syn181273)
    );
    X_BUF \syn20872/XUSED (
      .I (\syn20872/FROM ),
      .O (syn20872)
    );
    defparam C17641.INIT = 16'h8421;
    X_LUT4 C17641(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_minus1 [4]),
      .O (\syn182627/GROM )
    );
    X_BUF \syn182627/YUSED (
      .I (\syn182627/GROM ),
      .O (syn182627)
    );
    defparam C17617.INIT = 16'h8241;
    X_LUT4 C17617(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus3 [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [4]),
      .O (\syn182662/GROM )
    );
    defparam C17626.INIT = 16'h9009;
    X_LUT4 C17626(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_next [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [4]),
      .O (\syn182662/FROM )
    );
    X_BUF \syn182662/YUSED (
      .I (\syn182662/GROM ),
      .O (syn182679)
    );
    X_BUF \syn182662/XUSED (
      .I (\syn182662/FROM ),
      .O (syn182662)
    );
    defparam C19250.INIT = 16'hFFFB;
    X_LUT4 C19250(
      .ADR0 (syn19590),
      .ADR1 (syn19577),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_write_performed ),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .O (\bridge/pci_target_unit/fifos/pciw_rallow/GROM )
    );
    defparam C19251.INIT = 16'hE0C0;
    X_LUT4 C19251(
      .ADR0 (syn17011),
      .ADR1 (syn179021),
      .ADR2 (syn19577),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C983 ),
      .O (\bridge/pci_target_unit/fifos/pciw_rallow/FROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_rallow/YUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_rallow/GROM ),
      .O (\bridge/pci_target_unit/fifos/portB_enable )
    );
    X_BUF \bridge/pci_target_unit/fifos/pciw_rallow/XUSED (
      .I (\bridge/pci_target_unit/fifos/pciw_rallow/FROM ),
      .O (\bridge/pci_target_unit/fifos/pciw_rallow )
    );
    defparam C19170.INIT = 16'hF404;
    X_LUT4 C19170(
      .ADR0 (ADR_O[2]),
      .ADR1 (N_LED),
      .ADR2 (ADR_O[10]),
      .ADR3 (\CRT/wbs_pal_data [0]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[16]/GROM )
    );
    defparam C19219.INIT = 16'h00A0;
    X_LUT4 C19219(
      .ADR0 (\CRT/pix_start_addr [16]),
      .ADR1 (VCC),
      .ADR2 (ADR_O[2]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[16]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<16>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[16]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [0])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<16>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[16]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [16])
    );
    defparam C19162.INIT = 16'hF33F;
    X_LUT4 C19162(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_pci_am1_out [17]),
      .ADR2 (\bridge/conf_pci_ba1_out [17]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .O (\syn17052/GROM )
    );
    defparam C19856.INIT = 16'hC0C0;
    X_LUT4 C19856(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_pci_ba1_out [17]),
      .ADR2 (\bridge/conf_pci_am1_out [17]),
      .ADR3 (VCC),
      .O (\syn17052/FROM )
    );
    X_BUF \syn17052/YUSED (
      .I (\syn17052/GROM ),
      .O (syn19865)
    );
    X_BUF \syn17052/XUSED (
      .I (\syn17052/FROM ),
      .O (syn17052)
    );
    defparam C19066.INIT = 16'h5050;
    X_LUT4 C19066(
      .ADR0 (\CRT/drive_blank_reg ),
      .ADR1 (VCC),
      .ADR2 (\CRT/pal_pix_dat [5]),
      .ADR3 (VCC),
      .O (\rgb_int[4]/GROM )
    );
    defparam C19067.INIT = 16'h5050;
    X_LUT4 C19067(
      .ADR0 (\CRT/drive_blank_reg ),
      .ADR1 (VCC),
      .ADR2 (\CRT/pal_pix_dat [4]),
      .ADR3 (VCC),
      .O (\rgb_int[4]/FROM )
    );
    X_BUF \rgb_int<4>/YUSED (
      .I (\rgb_int[4]/GROM ),
      .O (rgb_int[5])
    );
    X_BUF \rgb_int<4>/XUSED (
      .I (\rgb_int[4]/FROM ),
      .O (rgb_int[4])
    );
    defparam C19058.INIT = 16'h00CC;
    X_LUT4 C19058(
      .ADR0 (VCC),
      .ADR1 (\CRT/pal_pix_dat [13]),
      .ADR2 (VCC),
      .ADR3 (\CRT/drive_blank_reg ),
      .O (\rgb_int[12]/GROM )
    );
    defparam C19059.INIT = 16'h3030;
    X_LUT4 C19059(
      .ADR0 (VCC),
      .ADR1 (\CRT/drive_blank_reg ),
      .ADR2 (\CRT/pal_pix_dat [12]),
      .ADR3 (VCC),
      .O (\rgb_int[12]/FROM )
    );
    X_BUF \rgb_int<12>/YUSED (
      .I (\rgb_int[12]/GROM ),
      .O (rgb_int[13])
    );
    X_BUF \rgb_int<12>/XUSED (
      .I (\rgb_int[12]/FROM ),
      .O (rgb_int[12])
    );
    defparam C18514.INIT = 16'hF888;
    X_LUT4 C18514(
      .ADR0 (\bridge/configuration/wb_err_data [17]),
      .ADR1 (\bridge/configuration/C1935 ),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/configuration/config_addr[17] ),
      .O (\syn180523/GROM )
    );
    defparam C18532.INIT = 16'hEAC0;
    X_LUT4 C18532(
      .ADR0 (\bridge/configuration/wb_err_data [16]),
      .ADR1 (\bridge/configuration/config_addr[16] ),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/configuration/C1935 ),
      .O (\syn180523/FROM )
    );
    X_BUF \syn180523/YUSED (
      .I (\syn180523/GROM ),
      .O (syn180564)
    );
    X_BUF \syn180523/XUSED (
      .I (\syn180523/FROM ),
      .O (syn180523)
    );
    defparam C18354.INIT = 16'hEAC0;
    X_LUT4 C18354(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [27]),
      .ADR1 (\bridge/conf_pci_am1_out [15]),
      .ADR2 (\bridge/configuration/C1989 ),
      .ADR3 (\bridge/configuration/C1987 ),
      .O (\syn180841/GROM )
    );
    defparam C18425.INIT = 16'hF888;
    X_LUT4 C18425(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [23]),
      .ADR1 (\bridge/configuration/C1989 ),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [23]),
      .ADR3 (\bridge/configuration/C1987 ),
      .O (\syn180841/FROM )
    );
    X_BUF \syn180841/YUSED (
      .I (\syn180841/GROM ),
      .O (syn181038)
    );
    X_BUF \syn180841/XUSED (
      .I (\syn180841/FROM ),
      .O (syn180841)
    );
    defparam C18346.INIT = 16'hECA0;
    X_LUT4 C18346(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [27]),
      .ADR1 (syn136384),
      .ADR2 (syn136386),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [27]),
      .O (\syn180957/GROM )
    );
    defparam C18382.INIT = 16'hF888;
    X_LUT4 C18382(
      .ADR0 (syn136384),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [25]),
      .ADR2 (syn136386),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [25]),
      .O (\syn180957/FROM )
    );
    X_BUF \syn180957/YUSED (
      .I (\syn180957/GROM ),
      .O (syn181058)
    );
    X_BUF \syn180957/XUSED (
      .I (\syn180957/FROM ),
      .O (syn180957)
    );
    defparam C18282.INIT = 16'hF888;
    X_LUT4 C18282(
      .ADR0 (\bridge/configuration/C2003 ),
      .ADR1 (\bridge/conf_pci_ba0_out [19]),
      .ADR2 (\bridge/configuration/C1925 ),
      .ADR3 (\bridge/configuration/icr_soft_res ),
      .O (\syn179985/GROM )
    );
    defparam C18722.INIT = 16'h8080;
    X_LUT4 C18722(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/configuration/serr_int_en ),
      .ADR2 (\bridge/configuration/C1925 ),
      .ADR3 (VCC),
      .O (\syn179985/FROM )
    );
    X_BUF \syn179985/YUSED (
      .I (\syn179985/GROM ),
      .O (syn181249)
    );
    X_BUF \syn179985/XUSED (
      .I (\syn179985/FROM ),
      .O (syn179985)
    );
    defparam C18274.INIT = 16'hECA0;
    X_LUT4 C18274(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [31]),
      .ADR1 (syn16931),
      .ADR2 (syn16919),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [31]),
      .O (\syn120400/GROM )
    );
    defparam C18293.INIT = 16'hECA0;
    X_LUT4 C18293(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [30]),
      .ADR1 (syn16919),
      .ADR2 (syn16931),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [30]),
      .O (\syn120400/FROM )
    );
    X_BUF \syn120400/YUSED (
      .I (\syn120400/GROM ),
      .O (syn120402)
    );
    X_BUF \syn120400/XUSED (
      .I (\syn120400/FROM ),
      .O (syn120400)
    );
    defparam C17802.INIT = 16'hFAFF;
    X_LUT4 C17802(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .ADR3 (syn17006),
      .O (\N12478/GROM )
    );
    defparam C17889.INIT = 16'hEEEA;
    X_LUT4 C17889(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .ADR1 (syn19713),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .O (\N12478/FROM )
    );
    X_BUF \N12478/YUSED (
      .I (\N12478/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C104/N6 )
    );
    X_BUF \N12478/XUSED (
      .I (\N12478/FROM ),
      .O (N12478)
    );
    defparam C17634.INIT = 16'h8241;
    X_LUT4 C17634(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_minus2 [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [3]),
      .O (\syn182610/GROM )
    );
    defparam C17653.INIT = 16'h9009;
    X_LUT4 C17653(
      .ADR0 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/rgrey_next [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pciw_fifo_ctrl/wgrey_addr [3]),
      .O (\syn182610/FROM )
    );
    X_BUF \syn182610/YUSED (
      .I (\syn182610/GROM ),
      .O (syn182650)
    );
    X_BUF \syn182610/XUSED (
      .I (\syn182610/FROM ),
      .O (syn182610)
    );
    defparam C19323.INIT = 16'h8421;
    X_LUT4 C19323(
      .ADR0 (\bridge/conf_pci_ba0_out [14]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .ADR3 (\bridge/conf_pci_ba0_out [13]),
      .O (\syn177733/GROM )
    );
    defparam C19812.INIT = 16'hF888;
    X_LUT4 C19812(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/pci_err_addr [26]),
      .ADR2 (\bridge/conf_pci_ba0_out [14]),
      .ADR3 (\bridge/configuration/C2370 ),
      .O (\syn177733/FROM )
    );
    X_BUF \syn177733/YUSED (
      .I (\syn177733/GROM ),
      .O (syn178850)
    );
    X_BUF \syn177733/XUSED (
      .I (\syn177733/FROM ),
      .O (syn177733)
    );
    defparam C19315.INIT = 16'h0001;
    X_LUT4 C19315(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/cnf_progress ),
      .ADR2 (\bridge/in_reg_irdy_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\syn16919/GROM )
    );
    X_BUF \syn16919/YUSED (
      .I (\syn16919/GROM ),
      .O (syn16919)
    );
    defparam C19171.INIT = 16'hF000;
    X_LUT4 C19171(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (ADR_O[10]),
      .ADR3 (\CRT/wbs_pal_data [1]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[17]/GROM )
    );
    defparam C19220.INIT = 16'h4400;
    X_LUT4 C19220(
      .ADR0 (ADR_O[10]),
      .ADR1 (ADR_O[2]),
      .ADR2 (VCC),
      .ADR3 (\CRT/pix_start_addr [17]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[17]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<17>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[17]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [1])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<17>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[17]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [17])
    );
    defparam C18515.INIT = 16'hEAC0;
    X_LUT4 C18515(
      .ADR0 (\bridge/configuration/C1989 ),
      .ADR1 (\bridge/configuration/pci_base_addr0 [17]),
      .ADR2 (\bridge/configuration/C2003 ),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [17]),
      .O (\syn180522/GROM )
    );
    defparam C18533.INIT = 16'hEAC0;
    X_LUT4 C18533(
      .ADR0 (\bridge/configuration/pci_base_addr0 [16]),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [16]),
      .ADR2 (\bridge/configuration/C1989 ),
      .ADR3 (\bridge/configuration/C2003 ),
      .O (\syn180522/FROM )
    );
    X_BUF \syn180522/YUSED (
      .I (\syn180522/GROM ),
      .O (syn180563)
    );
    X_BUF \syn180522/XUSED (
      .I (\syn180522/FROM ),
      .O (syn180522)
    );
    defparam C18451.INIT = 16'hF888;
    X_LUT4 C18451(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (\bridge/configuration/wb_err_data [21]),
      .ADR2 (\bridge/configuration/config_addr[21] ),
      .ADR3 (\bridge/configuration/C1929 ),
      .O (\syn180701/GROM )
    );
    defparam C18467.INIT = 16'hEAC0;
    X_LUT4 C18467(
      .ADR0 (\bridge/configuration/config_addr[20] ),
      .ADR1 (\bridge/configuration/C1935 ),
      .ADR2 (\bridge/configuration/wb_err_data [20]),
      .ADR3 (\bridge/configuration/C1929 ),
      .O (\syn180701/FROM )
    );
    X_BUF \syn180701/YUSED (
      .I (\syn180701/GROM ),
      .O (syn180747)
    );
    X_BUF \syn180701/XUSED (
      .I (\syn180701/FROM ),
      .O (syn180701)
    );
    defparam C18427.INIT = 16'hEA00;
    X_LUT4 C18427(
      .ADR0 (\bridge/configuration/C1953 ),
      .ADR1 (\bridge/configuration/wb_base_addr1 [23]),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [23]),
      .O (\syn21246/GROM )
    );
    defparam C18442.INIT = 16'hEA00;
    X_LUT4 C18442(
      .ADR0 (\bridge/configuration/C1953 ),
      .ADR1 (\bridge/configuration/wb_base_addr1 [22]),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [22]),
      .O (\syn21246/FROM )
    );
    X_BUF \syn21246/YUSED (
      .I (\syn21246/GROM ),
      .O (syn21285)
    );
    X_BUF \syn21246/XUSED (
      .I (\syn21246/FROM ),
      .O (syn21246)
    );
    defparam C18419.INIT = 16'h8C80;
    X_LUT4 C18419(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [23]),
      .ADR1 (syn19366),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [23]),
      .O (\syn180669/GROM )
    );
    defparam C18482.INIT = 16'hA0C0;
    X_LUT4 C18482(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [19]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [19]),
      .ADR2 (syn19366),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .O (\syn180669/FROM )
    );
    X_BUF \syn180669/YUSED (
      .I (\syn180669/GROM ),
      .O (syn180852)
    );
    X_BUF \syn180669/XUSED (
      .I (\syn180669/FROM ),
      .O (syn180669)
    );
    defparam C18283.INIT = 16'hFEFC;
    X_LUT4 C18283(
      .ADR0 (syn17049),
      .ADR1 (syn48754),
      .ADR2 (syn21610),
      .ADR3 (syn60110),
      .O (\bridge/configuration/C287/N3/GROM )
    );
    defparam C18826.INIT = 16'h4040;
    X_LUT4 C18826(
      .ADR0 (\bridge/in_reg_cbe_out [0]),
      .ADR1 (syn60110),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (VCC),
      .O (\bridge/configuration/C287/N3/FROM )
    );
    X_BUF \bridge/configuration/C287/N3/YUSED (
      .I (\bridge/configuration/C287/N3/GROM ),
      .O (syn181253)
    );
    X_BUF \bridge/configuration/C287/N3/XUSED (
      .I (\bridge/configuration/C287/N3/FROM ),
      .O (\bridge/configuration/C287/N3 )
    );
    defparam C19500.INIT = 16'hECA0;
    X_LUT4 C19500(
      .ADR0 (\bridge/conf_cache_line_size_out [1]),
      .ADR1 (\bridge/configuration/interrupt_line [1]),
      .ADR2 (syn17067),
      .ADR3 (syn17083),
      .O (\syn18659/GROM )
    );
    defparam C19560.INIT = 16'hA0A0;
    X_LUT4 C19560(
      .ADR0 (\bridge/conf_cache_line_size_out [7]),
      .ADR1 (VCC),
      .ADR2 (syn17067),
      .ADR3 (VCC),
      .O (\syn18659/FROM )
    );
    X_BUF \syn18659/YUSED (
      .I (\syn18659/GROM ),
      .O (syn178495)
    );
    X_BUF \syn18659/XUSED (
      .I (\syn18659/FROM ),
      .O (syn18659)
    );
    defparam C19404.INIT = 16'h555F;
    X_LUT4 C19404(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/write_req_int ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_rdy_out ),
      .O (\syn16939/GROM )
    );
    defparam C19470.INIT = 16'h0800;
    X_LUT4 C19470(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_rdy_out ),
      .ADR1 (syn17023),
      .ADR2 (N12594),
      .ADR3 (N12359),
      .O (\syn16939/FROM )
    );
    X_BUF \syn16939/YUSED (
      .I (\syn16939/GROM ),
      .O (syn178714)
    );
    X_BUF \syn16939/XUSED (
      .I (\syn16939/FROM ),
      .O (syn16939)
    );
    defparam C19324.INIT = 16'h8484;
    X_LUT4 C19324(
      .ADR0 (\bridge/conf_pci_ba0_out [18]),
      .ADR1 (\bridge/conf_mem_space_enable_out ),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .ADR3 (VCC),
      .O (\syn17875/GROM )
    );
    defparam C19889.INIT = 16'h8888;
    X_LUT4 C19889(
      .ADR0 (syn16930),
      .ADR1 (\bridge/conf_pci_ba0_out [18]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn17875/FROM )
    );
    X_BUF \syn17875/YUSED (
      .I (\syn17875/GROM ),
      .O (syn178847)
    );
    X_BUF \syn17875/XUSED (
      .I (\syn17875/FROM ),
      .O (syn17875)
    );
    defparam C19180.INIT = 16'hEC20;
    X_LUT4 C19180(
      .ADR0 (\CRT/pix_start_addr [10]),
      .ADR1 (ADR_O[10]),
      .ADR2 (ADR_O[2]),
      .ADR3 (\CRT/wbs_pal_data [10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[26]/GROM )
    );
    defparam C19229.INIT = 16'h5000;
    X_LUT4 C19229(
      .ADR0 (ADR_O[10]),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [26]),
      .ADR3 (ADR_O[2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[26]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<26>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[26]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [10])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<26>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[26]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [26])
    );
    defparam C19172.INIT = 16'hF808;
    X_LUT4 C19172(
      .ADR0 (ADR_O[2]),
      .ADR1 (\CRT/pix_start_addr [2]),
      .ADR2 (ADR_O[10]),
      .ADR3 (\CRT/wbs_pal_data [2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[18]/GROM )
    );
    defparam C19221.INIT = 16'h0A00;
    X_LUT4 C19221(
      .ADR0 (ADR_O[2]),
      .ADR1 (VCC),
      .ADR2 (ADR_O[10]),
      .ADR3 (\CRT/pix_start_addr [18]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[18]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<18>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[18]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [2])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<18>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[18]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [18])
    );
    defparam C18516.INIT = 16'hEAC0;
    X_LUT4 C18516(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (\bridge/configuration/C1987 ),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [17]),
      .ADR3 (\bridge/configuration/wb_tran_addr1 [17]),
      .O (\syn180521/GROM )
    );
    defparam C18534.INIT = 16'hECA0;
    X_LUT4 C18534(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (\bridge/configuration/C1987 ),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [16]),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [16]),
      .O (\syn180521/FROM )
    );
    X_BUF \syn180521/YUSED (
      .I (\syn180521/GROM ),
      .O (syn180562)
    );
    X_BUF \syn180521/XUSED (
      .I (\syn180521/FROM ),
      .O (syn180521)
    );
    defparam C18452.INIT = 16'hF888;
    X_LUT4 C18452(
      .ADR0 (\bridge/configuration/pci_addr_mask1 [21]),
      .ADR1 (\bridge/configuration/C1989 ),
      .ADR2 (\bridge/configuration/C2003 ),
      .ADR3 (\bridge/configuration/pci_base_addr0 [21]),
      .O (\syn180700/GROM )
    );
    defparam C18468.INIT = 16'hF888;
    X_LUT4 C18468(
      .ADR0 (\bridge/configuration/pci_base_addr0 [20]),
      .ADR1 (\bridge/configuration/C2003 ),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [20]),
      .ADR3 (\bridge/configuration/C1989 ),
      .O (\syn180700/FROM )
    );
    X_BUF \syn180700/YUSED (
      .I (\syn180700/GROM ),
      .O (syn180746)
    );
    X_BUF \syn180700/XUSED (
      .I (\syn180700/FROM ),
      .O (syn180700)
    );
    defparam C18372.INIT = 16'hF888;
    X_LUT4 C18372(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [26]),
      .ADR1 (\bridge/configuration/C1951 ),
      .ADR2 (syn60110),
      .ADR3 (syn17055),
      .O (\syn180840/GROM )
    );
    defparam C18426.INIT = 16'hF888;
    X_LUT4 C18426(
      .ADR0 (syn17058),
      .ADR1 (syn60110),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [23]),
      .ADR3 (\bridge/configuration/C1951 ),
      .O (\syn180840/FROM )
    );
    X_BUF \syn180840/YUSED (
      .I (\syn180840/GROM ),
      .O (syn180992)
    );
    X_BUF \syn180840/XUSED (
      .I (\syn180840/FROM ),
      .O (syn180840)
    );
    defparam C18364.INIT = 16'hECA0;
    X_LUT4 C18364(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [26]),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [26]),
      .O (\syn180951/GROM )
    );
    defparam C18385.INIT = 16'hECA0;
    X_LUT4 C18385(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [25]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_data_out [25]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (syn20493),
      .O (\syn180951/FROM )
    );
    X_BUF \syn180951/YUSED (
      .I (\syn180951/GROM ),
      .O (syn180971)
    );
    X_BUF \syn180951/XUSED (
      .I (\syn180951/FROM ),
      .O (syn180951)
    );
    defparam C18356.INIT = 16'hE0C0;
    X_LUT4 C18356(
      .ADR0 (\bridge/conf_wb_ba1_out [15]),
      .ADR1 (\bridge/configuration/C1953 ),
      .ADR2 (\bridge/conf_wb_am1_out [15]),
      .ADR3 (\bridge/configuration/C1955 ),
      .O (\syn17971/GROM )
    );
    defparam C19832.INIT = 16'hC8C0;
    X_LUT4 C19832(
      .ADR0 (\bridge/conf_wb_ba1_out [15]),
      .ADR1 (\bridge/conf_wb_am1_out [15]),
      .ADR2 (\bridge/configuration/C2320 ),
      .ADR3 (\bridge/configuration/C2322 ),
      .O (\syn17971/FROM )
    );
    X_BUF \syn17971/YUSED (
      .I (\syn17971/GROM ),
      .O (syn21448)
    );
    X_BUF \syn17971/XUSED (
      .I (\syn17971/FROM ),
      .O (syn17971)
    );
    defparam C18292.INIT = 16'hE0A0;
    X_LUT4 C18292(
      .ADR0 (syn120400),
      .ADR1 (\bridge/conf_pci_ba0_out [18]),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn16929),
      .O (\syn181166/GROM )
    );
    defparam C18309.INIT = 16'hA888;
    X_LUT4 C18309(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn120398),
      .ADR2 (\bridge/conf_pci_ba0_out [17]),
      .ADR3 (syn16929),
      .O (\syn181166/FROM )
    );
    X_BUF \syn181166/YUSED (
      .I (\syn181166/GROM ),
      .O (syn181218)
    );
    X_BUF \syn181166/XUSED (
      .I (\syn181166/FROM ),
      .O (syn181166)
    );
    defparam C18284.INIT = 16'hC000;
    X_LUT4 C18284(
      .ADR0 (VCC),
      .ADR1 (\bridge/conf_wb_am1_out [19]),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/conf_wb_ba1_out [19]),
      .O (\syn177524/GROM )
    );
    defparam C19903.INIT = 16'h8800;
    X_LUT4 C19903(
      .ADR0 (syn16917),
      .ADR1 (\bridge/conf_wb_am1_out [19]),
      .ADR2 (VCC),
      .ADR3 (syn24500),
      .O (\syn177524/FROM )
    );
    X_BUF \syn177524/YUSED (
      .I (\syn177524/GROM ),
      .O (syn21610)
    );
    X_BUF \syn177524/XUSED (
      .I (\syn177524/FROM ),
      .O (syn177524)
    );
    defparam C17812.INIT = 16'hFFF0;
    X_LUT4 C17812(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn23069),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/reset_rty_cnt ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en/GROM )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/rty_cnt_clk_en )
    );
    defparam C19501.INIT = 16'hECA0;
    X_LUT4 C19501(
      .ADR0 (syn24559),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [1]),
      .ADR2 (\bridge/conf_mem_space_enable_out ),
      .ADR3 (syn17745),
      .O (\syn177830/GROM )
    );
    defparam C19778.INIT = 16'hEAC0;
    X_LUT4 C19778(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [24]),
      .ADR1 (\bridge/configuration/status_bit8 ),
      .ADR2 (syn24559),
      .ADR3 (syn17745),
      .O (\syn177830/FROM )
    );
    X_BUF \syn177830/YUSED (
      .I (\syn177830/GROM ),
      .O (syn178494)
    );
    X_BUF \syn177830/XUSED (
      .I (\syn177830/FROM ),
      .O (syn177830)
    );
    defparam C19325.INIT = 16'h8421;
    X_LUT4 C19325(
      .ADR0 (\bridge/conf_pci_ba0_out [16]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .ADR3 (\bridge/conf_pci_ba0_out [15]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[28]/GROM )
    );
    defparam C19381.INIT = 16'hFFAA;
    X_LUT4 C19381(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[28]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<28>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[28]/GROM ),
      .O (syn178849)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<28>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[28]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [28])
    );
    defparam C19181.INIT = 16'hCAC0;
    X_LUT4 C19181(
      .ADR0 (ADR_O[2]),
      .ADR1 (\CRT/wbs_pal_data [11]),
      .ADR2 (ADR_O[10]),
      .ADR3 (\CRT/pix_start_addr [11]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[27]/GROM )
    );
    defparam C19230.INIT = 16'h4400;
    X_LUT4 C19230(
      .ADR0 (ADR_O[10]),
      .ADR1 (\CRT/pix_start_addr [27]),
      .ADR2 (VCC),
      .ADR3 (ADR_O[2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[27]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<27>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[27]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [11])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<27>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[27]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [27])
    );
    defparam C19173.INIT = 16'hACA0;
    X_LUT4 C19173(
      .ADR0 (\CRT/wbs_pal_data [3]),
      .ADR1 (\CRT/pix_start_addr [3]),
      .ADR2 (ADR_O[10]),
      .ADR3 (ADR_O[2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[19]/GROM )
    );
    defparam C19222.INIT = 16'h00A0;
    X_LUT4 C19222(
      .ADR0 (ADR_O[2]),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [19]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[19]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<19>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[19]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [3])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<19>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[19]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [19])
    );
    defparam C18453.INIT = 16'hECA0;
    X_LUT4 C18453(
      .ADR0 (\bridge/configuration/C1987 ),
      .ADR1 (\bridge/configuration/C1951 ),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [21]),
      .ADR3 (\bridge/configuration/wb_tran_addr1 [21]),
      .O (\syn180699/GROM )
    );
    defparam C18469.INIT = 16'hEAC0;
    X_LUT4 C18469(
      .ADR0 (\bridge/configuration/C1987 ),
      .ADR1 (\bridge/configuration/C1951 ),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [20]),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [20]),
      .O (\syn180699/FROM )
    );
    X_BUF \syn180699/YUSED (
      .I (\syn180699/GROM ),
      .O (syn180745)
    );
    X_BUF \syn180699/XUSED (
      .I (\syn180699/FROM ),
      .O (syn180699)
    );
    defparam C18285.INIT = 16'hECA0;
    X_LUT4 C18285(
      .ADR0 (\bridge/configuration/C1989 ),
      .ADR1 (\bridge/configuration/C1987 ),
      .ADR2 (\bridge/conf_pci_am1_out [19]),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [31]),
      .O (\syn181194/GROM )
    );
    defparam C18298.INIT = 16'hEAC0;
    X_LUT4 C18298(
      .ADR0 (\bridge/configuration/C1989 ),
      .ADR1 (\bridge/configuration/C1987 ),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [30]),
      .ADR3 (\bridge/conf_pci_am1_out [18]),
      .O (\syn181194/FROM )
    );
    X_BUF \syn181194/YUSED (
      .I (\syn181194/GROM ),
      .O (syn181248)
    );
    X_BUF \syn181194/XUSED (
      .I (\syn181194/FROM ),
      .O (syn181194)
    );
    defparam C17725.INIT = 16'hFFCF;
    X_LUT4 C17725(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync_comp_flush_out ),
      .ADR2 (N_RST),
      .ADR3 (\bridge/wishbone_slave_unit/wbs_sm_wbr_flush_out ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear/GROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear/GROM ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear )
    );
    defparam C19318.INIT = 16'h222E;
    X_LUT4 C19318(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/N5157 ),
      .ADR1 (\bridge/in_reg_cbe_out [3]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/conf_addr_out [0]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/conf_addr_out [1]),
      .O (\bridge/pci_target_unit/pci_target_sm/cnf_progress/GROM )
    );
    defparam C19169.INIT = 16'h2000;
    X_LUT4 C19169(
      .ADR0 (\bridge/in_reg_idsel_out ),
      .ADR1 (\bridge/in_reg_cbe_out [2]),
      .ADR2 (\bridge/in_reg_cbe_out [3]),
      .ADR3 (\bridge/in_reg_cbe_out [1]),
      .O (\bridge/pci_target_unit/pci_target_sm/cnf_progress/FROM )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/cnf_progress/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/cnf_progress/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/cnf_progress/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/cnf_progress/GROM ),
      .O (syn19380)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/cnf_progress/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/cnf_progress/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/config_access )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/cnf_progress_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/cnf_progress/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/cnf_progress/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/cnf_progress )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/cnf_progress/FFX/ASYNC_FF_GSR_OR_144 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/cnf_progress/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/cnf_progress/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19270.INIT = 16'hBB88;
    X_LUT4 C19270(
      .ADR0 (\bridge/pci_target_unit/pcit_if_addr_out [21]),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[22]/GROM )
    );
    defparam C19271.INIT = 16'hF3C0;
    X_LUT4 C19271(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR2 (\bridge/pci_target_unit/pcit_if_addr_out [22]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[22]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<22>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[22]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [21])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<22>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[22]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [22])
    );
    defparam C19190.INIT = 16'hCACA;
    X_LUT4 C19190(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [4]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[4]/GROM )
    );
    defparam C19333.INIT = 16'hFFAA;
    X_LUT4 C19333(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[4]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<4>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[4]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [4])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<4>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[4]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [4])
    );
    defparam C19182.INIT = 16'hF808;
    X_LUT4 C19182(
      .ADR0 (\CRT/pix_start_addr [12]),
      .ADR1 (ADR_O[2]),
      .ADR2 (ADR_O[10]),
      .ADR3 (\CRT/wbs_pal_data [12]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[28]/GROM )
    );
    defparam C19231.INIT = 16'h0088;
    X_LUT4 C19231(
      .ADR0 (ADR_O[2]),
      .ADR1 (\CRT/pix_start_addr [28]),
      .ADR2 (VCC),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[28]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<28>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[28]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [12])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<28>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[28]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [28])
    );
    defparam C19174.INIT = 16'hCCA0;
    X_LUT4 C19174(
      .ADR0 (\CRT/pix_start_addr [4]),
      .ADR1 (\CRT/wbs_pal_data [4]),
      .ADR2 (ADR_O[2]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[20]/GROM )
    );
    defparam C19223.INIT = 16'h0A00;
    X_LUT4 C19223(
      .ADR0 (\CRT/pix_start_addr [20]),
      .ADR1 (VCC),
      .ADR2 (ADR_O[10]),
      .ADR3 (ADR_O[2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[20]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<20>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[20]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [4])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<20>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[20]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [20])
    );
    defparam C18630.INIT = 16'hF888;
    X_LUT4 C18630(
      .ADR0 (syn17016),
      .ADR1 (\bridge/configuration/config_addr[10] ),
      .ADR2 (\bridge/conf_latency_tim_out [2]),
      .ADR3 (syn17102),
      .O (\syn180205/GROM )
    );
    defparam C18645.INIT = 16'hF888;
    X_LUT4 C18645(
      .ADR0 (syn17016),
      .ADR1 (\bridge/configuration/config_addr[9] ),
      .ADR2 (syn17102),
      .ADR3 (\bridge/conf_latency_tim_out [1]),
      .O (\syn180205/FROM )
    );
    X_BUF \syn180205/YUSED (
      .I (\syn180205/GROM ),
      .O (syn180244)
    );
    X_BUF \syn180205/XUSED (
      .I (\syn180205/FROM ),
      .O (syn180205)
    );
    defparam C18438.INIT = 16'hEAC0;
    X_LUT4 C18438(
      .ADR0 (\bridge/configuration/wb_err_addr [22]),
      .ADR1 (\bridge/configuration/C1935 ),
      .ADR2 (\bridge/configuration/wb_err_data [22]),
      .ADR3 (\bridge/configuration/C1937 ),
      .O (\syn180660/GROM )
    );
    defparam C18486.INIT = 16'hF888;
    X_LUT4 C18486(
      .ADR0 (\bridge/configuration/wb_err_addr [19]),
      .ADR1 (\bridge/configuration/C1937 ),
      .ADR2 (\bridge/configuration/wb_err_data [19]),
      .ADR3 (\bridge/configuration/C1935 ),
      .O (\syn180660/FROM )
    );
    X_BUF \syn180660/YUSED (
      .I (\syn180660/GROM ),
      .O (syn180793)
    );
    X_BUF \syn180660/XUSED (
      .I (\syn180660/FROM ),
      .O (syn180660)
    );
    defparam C18286.INIT = 16'hECA0;
    X_LUT4 C18286(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (\bridge/configuration/C1953 ),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [31]),
      .ADR3 (\bridge/conf_wb_am1_out [19]),
      .O (\syn21571/GROM )
    );
    defparam C18300.INIT = 16'hC8C0;
    X_LUT4 C18300(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/conf_wb_am1_out [18]),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/conf_wb_ba1_out [18]),
      .O (\syn21571/FROM )
    );
    X_BUF \syn21571/YUSED (
      .I (\syn21571/GROM ),
      .O (syn181247)
    );
    X_BUF \syn21571/XUSED (
      .I (\syn21571/FROM ),
      .O (syn21571)
    );
    defparam C19335.INIT = 16'hFFCC;
    X_LUT4 C19335(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[12]/GROM )
    );
    defparam C19341.INIT = 16'hFFCC;
    X_LUT4 C19341(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[12]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<12>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[12]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [6])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<12>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[12]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [12])
    );
    defparam C19263.INIT = 16'h8000;
    X_LUT4 C19263(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/rty_counter [3]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/rty_counter [1]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/rty_counter [0]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/rty_counter [2]),
      .O (\syn178999/GROM )
    );
    X_BUF \syn178999/YUSED (
      .I (\syn178999/GROM ),
      .O (syn178999)
    );
    defparam C19191.INIT = 16'hF3C0;
    X_LUT4 C19191(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR2 (\bridge/pci_target_unit/pcit_if_addr_out [5]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[6]/GROM )
    );
    defparam C19192.INIT = 16'hAACC;
    X_LUT4 C19192(
      .ADR0 (\bridge/pci_target_unit/pcit_if_addr_out [6]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[6]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<6>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[6]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [5])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<6>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[6]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [6])
    );
    defparam C19183.INIT = 16'hAAC0;
    X_LUT4 C19183(
      .ADR0 (\CRT/wbs_pal_data [13]),
      .ADR1 (\CRT/pix_start_addr [13]),
      .ADR2 (ADR_O[2]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[29]/GROM )
    );
    defparam C19232.INIT = 16'h0C00;
    X_LUT4 C19232(
      .ADR0 (VCC),
      .ADR1 (\CRT/pix_start_addr [29]),
      .ADR2 (ADR_O[10]),
      .ADR3 (ADR_O[2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[29]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<29>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[29]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [13])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<29>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[29]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [29])
    );
    defparam C19175.INIT = 16'hB888;
    X_LUT4 C19175(
      .ADR0 (\CRT/wbs_pal_data [5]),
      .ADR1 (ADR_O[10]),
      .ADR2 (ADR_O[2]),
      .ADR3 (\CRT/pix_start_addr [5]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[21]/GROM )
    );
    defparam C19224.INIT = 16'h4040;
    X_LUT4 C19224(
      .ADR0 (ADR_O[10]),
      .ADR1 (\CRT/pix_start_addr [21]),
      .ADR2 (ADR_O[2]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[21]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<21>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[21]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [5])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<21>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[21]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [21])
    );
    defparam C18703.INIT = 16'hEAC0;
    X_LUT4 C18703(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [4]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [4]),
      .ADR3 (syn20493),
      .O (\syn179931/GROM )
    );
    defparam C18739.INIT = 16'hECA0;
    X_LUT4 C18739(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [2]),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_data_out [2]),
      .O (\syn179931/FROM )
    );
    X_BUF \syn179931/YUSED (
      .I (\syn179931/GROM ),
      .O (syn180012)
    );
    X_BUF \syn179931/XUSED (
      .I (\syn179931/FROM ),
      .O (syn179931)
    );
    defparam C18631.INIT = 16'hC000;
    X_LUT4 C18631(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/C1973 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/configuration/pci_error_rty_exp_set ),
      .O (\syn180138/GROM )
    );
    defparam C18658.INIT = 16'h8000;
    X_LUT4 C18658(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/conf_pci_err_pending_out ),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (\bridge/configuration/C1973 ),
      .O (\syn180138/FROM )
    );
    X_BUF \syn180138/YUSED (
      .I (\syn180138/GROM ),
      .O (syn20796)
    );
    X_BUF \syn180138/XUSED (
      .I (\syn180138/FROM ),
      .O (syn180138)
    );
    defparam C18543.INIT = 16'hAA80;
    X_LUT4 C18543(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn16927),
      .ADR2 (syn17066),
      .ADR3 (syn120386),
      .O (\syn20484/GROM )
    );
    defparam C18774.INIT = 16'h8800;
    X_LUT4 C18774(
      .ADR0 (\bridge/conf_pci_mem_io1_out ),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (VCC),
      .ADR3 (syn16927),
      .O (\syn20484/FROM )
    );
    X_BUF \syn20484/YUSED (
      .I (\syn20484/GROM ),
      .O (syn180489)
    );
    X_BUF \syn20484/XUSED (
      .I (\syn20484/FROM ),
      .O (syn20484)
    );
    defparam C18519.INIT = 16'hA8A0;
    X_LUT4 C18519(
      .ADR0 (\bridge/configuration/wb_addr_mask1 [17]),
      .ADR1 (\bridge/configuration/wb_base_addr1 [17]),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/configuration/C1955 ),
      .O (\syn178054/GROM )
    );
    defparam C19693.INIT = 16'hF8F0;
    X_LUT4 C19693(
      .ADR0 (\bridge/configuration/wb_addr_mask1 [17]),
      .ADR1 (\bridge/configuration/wb_base_addr1 [17]),
      .ADR2 (\bridge/configuration/C2368 ),
      .ADR3 (\bridge/configuration/C2322 ),
      .O (\syn178054/FROM )
    );
    X_BUF \syn178054/YUSED (
      .I (\syn178054/GROM ),
      .O (syn21053)
    );
    X_BUF \syn178054/XUSED (
      .I (\syn178054/FROM ),
      .O (syn178054)
    );
    defparam C18391.INIT = 16'hF888;
    X_LUT4 C18391(
      .ADR0 (\bridge/conf_pci_am1_out [13]),
      .ADR1 (\bridge/configuration/C1989 ),
      .ADR2 (\bridge/conf_pci_ba0_out [13]),
      .ADR3 (\bridge/configuration/C2003 ),
      .O (\syn180884/GROM )
    );
    defparam C18408.INIT = 16'hECA0;
    X_LUT4 C18408(
      .ADR0 (\bridge/configuration/C2003 ),
      .ADR1 (\bridge/configuration/C1989 ),
      .ADR2 (\bridge/conf_pci_ba0_out [12]),
      .ADR3 (\bridge/conf_pci_am1_out [12]),
      .O (\syn180884/FROM )
    );
    X_BUF \syn180884/YUSED (
      .I (\syn180884/GROM ),
      .O (syn180936)
    );
    X_BUF \syn180884/XUSED (
      .I (\syn180884/FROM ),
      .O (syn180884)
    );
    defparam C18383.INIT = 16'hEA00;
    X_LUT4 C18383(
      .ADR0 (syn17104),
      .ADR1 (syn16929),
      .ADR2 (\bridge/conf_pci_ba0_out [13]),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn180907/GROM )
    );
    defparam C18397.INIT = 16'hF080;
    X_LUT4 C18397(
      .ADR0 (\bridge/conf_pci_ba0_out [12]),
      .ADR1 (syn16929),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn120394),
      .O (\syn180907/FROM )
    );
    X_BUF \syn180907/YUSED (
      .I (\syn180907/GROM ),
      .O (syn180960)
    );
    X_BUF \syn180907/XUSED (
      .I (\syn180907/FROM ),
      .O (syn180907)
    );
    defparam C18279.INIT = 16'hEAC0;
    X_LUT4 C18279(
      .ADR0 (\bridge/configuration/C1973 ),
      .ADR1 (\bridge/configuration/pci_err_addr [31]),
      .ADR2 (\bridge/configuration/C1971 ),
      .ADR3 (\bridge/configuration/pci_err_cs_bit31_24 [31]),
      .O (\syn181146/GROM )
    );
    defparam C18317.INIT = 16'hEAC0;
    X_LUT4 C18317(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/configuration/C1973 ),
      .ADR2 (\bridge/configuration/pci_err_cs_bit31_24 [29]),
      .ADR3 (\bridge/configuration/pci_err_addr [29]),
      .O (\syn181146/FROM )
    );
    X_BUF \syn181146/YUSED (
      .I (\syn181146/GROM ),
      .O (syn181252)
    );
    X_BUF \syn181146/XUSED (
      .I (\syn181146/FROM ),
      .O (syn181146)
    );
    defparam C18199.INIT = 16'h6FF6;
    X_LUT4 C18199(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/inGreyCount [1]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/outGreyCount [1]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/inGreyCount [0]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/outGreyCount [0]),
      .O (\syn181403/GROM )
    );
    X_BUF \syn181403/YUSED (
      .I (\syn181403/GROM ),
      .O (syn181403)
    );
    defparam C17719.INIT = 16'h9009;
    X_LUT4 C17719(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [3]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_next [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [2]),
      .O (\syn182474/GROM )
    );
    defparam C17723.INIT = 16'h6FF6;
    X_LUT4 C17723(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [3]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rgrey_addr [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [2]),
      .O (\syn182474/FROM )
    );
    X_BUF \syn182474/YUSED (
      .I (\syn182474/GROM ),
      .O (syn182485)
    );
    X_BUF \syn182474/XUSED (
      .I (\syn182474/FROM ),
      .O (syn182474)
    );
    defparam C19600.INIT = 16'h8888;
    X_LUT4 C19600(
      .ADR0 (\bridge/configuration/C2334 ),
      .ADR1 (syn16917),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn17073/GROM )
    );
    defparam C19603.INIT = 16'hCC00;
    X_LUT4 C19603(
      .ADR0 (VCC),
      .ADR1 (syn16917),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn17073/FROM )
    );
    X_BUF \syn17073/YUSED (
      .I (\syn17073/GROM ),
      .O (syn17072)
    );
    X_BUF \syn17073/XUSED (
      .I (\syn17073/FROM ),
      .O (syn17073)
    );
    defparam C19520.INIT = 16'h8800;
    X_LUT4 C19520(
      .ADR0 (syn177632),
      .ADR1 (\bridge/configuration/pci_img_ctrl1 [2]),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C3488 ),
      .O (\syn18756/GROM )
    );
    X_BUF \syn18756/YUSED (
      .I (\syn18756/GROM ),
      .O (syn18756)
    );
    defparam C19280.INIT = 16'hEE22;
    X_LUT4 C19280(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pcit_if_addr_out [31]),
      .O (\syn178848/GROM )
    );
    defparam C19326.INIT = 16'h8241;
    X_LUT4 C19326(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .ADR2 (\bridge/conf_pci_ba0_out [17]),
      .ADR3 (\bridge/conf_pci_ba0_out [19]),
      .O (\syn178848/FROM )
    );
    X_BUF \syn178848/YUSED (
      .I (\syn178848/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [31])
    );
    X_BUF \syn178848/XUSED (
      .I (\syn178848/FROM ),
      .O (syn178848)
    );
    defparam C19272.INIT = 16'hF0AA;
    X_LUT4 C19272(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pcit_if_addr_out [23]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[24]/GROM )
    );
    defparam C19273.INIT = 16'hAACC;
    X_LUT4 C19273(
      .ADR0 (\bridge/pci_target_unit/pcit_if_addr_out [24]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[24]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<24>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[24]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [23])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<24>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[24]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [24])
    );
    defparam C19264.INIT = 16'h8000;
    X_LUT4 C19264(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/rty_counter [7]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/rty_counter [6]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/rty_counter [4]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/rty_counter [5]),
      .O (\syn178998/GROM )
    );
    X_BUF \syn178998/YUSED (
      .I (\syn178998/GROM ),
      .O (syn178998)
    );
    defparam C19184.INIT = 16'hE4A0;
    X_LUT4 C19184(
      .ADR0 (ADR_O[10]),
      .ADR1 (ADR_O[2]),
      .ADR2 (\CRT/wbs_pal_data [14]),
      .ADR3 (\CRT/pix_start_addr [14]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[30]/GROM )
    );
    defparam C19233.INIT = 16'h2200;
    X_LUT4 C19233(
      .ADR0 (\CRT/pix_start_addr [30]),
      .ADR1 (ADR_O[10]),
      .ADR2 (VCC),
      .ADR3 (ADR_O[2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[30]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<30>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[30]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [14])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<30>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[30]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [30])
    );
    defparam C19176.INIT = 16'hF088;
    X_LUT4 C19176(
      .ADR0 (ADR_O[2]),
      .ADR1 (\CRT/pix_start_addr [6]),
      .ADR2 (\CRT/wbs_pal_data [6]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[22]/GROM )
    );
    defparam C19225.INIT = 16'h2200;
    X_LUT4 C19225(
      .ADR0 (ADR_O[2]),
      .ADR1 (ADR_O[10]),
      .ADR2 (VCC),
      .ADR3 (\CRT/pix_start_addr [22]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[22]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<22>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[22]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [6])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<22>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[22]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [22])
    );
    defparam C18608.INIT = 16'hC8C0;
    X_LUT4 C18608(
      .ADR0 (\bridge/configuration/wb_base_addr1 [12]),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [12]),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/configuration/C1955 ),
      .O (\syn178236/GROM )
    );
    defparam C19621.INIT = 16'hEAAA;
    X_LUT4 C19621(
      .ADR0 (\bridge/configuration/C2368 ),
      .ADR1 (\bridge/configuration/wb_base_addr1 [12]),
      .ADR2 (\bridge/configuration/C2322 ),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [12]),
      .O (\syn178236/FROM )
    );
    X_BUF \syn178236/YUSED (
      .I (\syn178236/GROM ),
      .O (syn20853)
    );
    X_BUF \syn178236/XUSED (
      .I (\syn178236/FROM ),
      .O (syn178236)
    );
    defparam C18560.INIT = 16'hF800;
    X_LUT4 C18560(
      .ADR0 (syn17068),
      .ADR1 (syn16927),
      .ADR2 (syn120384),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn20909/GROM )
    );
    defparam C18577.INIT = 16'h8000;
    X_LUT4 C18577(
      .ADR0 (\bridge/configuration/pci_base_addr1 [13]),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [13]),
      .ADR2 (syn16927),
      .ADR3 (\bridge/out_bckp_tar_ad_en_out ),
      .O (\syn20909/FROM )
    );
    X_BUF \syn20909/YUSED (
      .I (\syn20909/GROM ),
      .O (syn180439)
    );
    X_BUF \syn20909/XUSED (
      .I (\syn20909/FROM ),
      .O (syn20909)
    );
    defparam C18552.INIT = 16'hCC80;
    X_LUT4 C18552(
      .ADR0 (\bridge/configuration/wb_base_addr1 [15]),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [15]),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/configuration/C1953 ),
      .O (\syn20934/GROM )
    );
    defparam C18570.INIT = 16'hEA00;
    X_LUT4 C18570(
      .ADR0 (\bridge/configuration/C1953 ),
      .ADR1 (\bridge/configuration/wb_base_addr1 [14]),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [14]),
      .O (\syn20934/FROM )
    );
    X_BUF \syn20934/YUSED (
      .I (\syn20934/GROM ),
      .O (syn20974)
    );
    X_BUF \syn20934/XUSED (
      .I (\syn20934/FROM ),
      .O (syn20934)
    );
    defparam C18472.INIT = 16'hA888;
    X_LUT4 C18472(
      .ADR0 (\bridge/configuration/wb_addr_mask1 [20]),
      .ADR1 (\bridge/configuration/C1953 ),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/configuration/wb_base_addr1 [20]),
      .O (\syn177954/GROM )
    );
    defparam C19732.INIT = 16'hEAAA;
    X_LUT4 C19732(
      .ADR0 (\bridge/configuration/C2368 ),
      .ADR1 (\bridge/configuration/C2322 ),
      .ADR2 (\bridge/configuration/wb_base_addr1 [20]),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [20]),
      .O (\syn177954/FROM )
    );
    X_BUF \syn177954/YUSED (
      .I (\syn177954/GROM ),
      .O (syn21170)
    );
    X_BUF \syn177954/XUSED (
      .I (\syn177954/FROM ),
      .O (syn177954)
    );
    defparam C18464.INIT = 16'hEAC0;
    X_LUT4 C18464(
      .ADR0 (syn136384),
      .ADR1 (syn136386),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [20]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [20]),
      .O (\syn180626/GROM )
    );
    defparam C18495.INIT = 16'hECA0;
    X_LUT4 C18495(
      .ADR0 (syn136384),
      .ADR1 (syn136386),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [18]),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [18]),
      .O (\syn180626/FROM )
    );
    X_BUF \syn180626/YUSED (
      .I (\syn180626/GROM ),
      .O (syn180717)
    );
    X_BUF \syn180626/XUSED (
      .I (\syn180626/FROM ),
      .O (syn180626)
    );
    defparam C18456.INIT = 16'hF800;
    X_LUT4 C18456(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/configuration/wb_base_addr1 [21]),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [21]),
      .O (\syn177921/GROM )
    );
    defparam C19745.INIT = 16'hEAAA;
    X_LUT4 C19745(
      .ADR0 (\bridge/configuration/C2368 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [21]),
      .ADR2 (\bridge/configuration/wb_base_addr1 [21]),
      .ADR3 (\bridge/configuration/C2322 ),
      .O (\syn177921/FROM )
    );
    X_BUF \syn177921/YUSED (
      .I (\syn177921/GROM ),
      .O (syn21208)
    );
    X_BUF \syn177921/XUSED (
      .I (\syn177921/FROM ),
      .O (syn177921)
    );
    defparam C18376.INIT = 16'hECA0;
    X_LUT4 C18376(
      .ADR0 (\bridge/configuration/C1941 ),
      .ADR1 (\bridge/configuration/wb_err_addr [26]),
      .ADR2 (\bridge/configuration/wb_err_cs_bit31_24 [26]),
      .ADR3 (\bridge/configuration/C1937 ),
      .O (\syn179848/GROM )
    );
    defparam C18791.INIT = 16'hECA0;
    X_LUT4 C18791(
      .ADR0 (\bridge/configuration/C1937 ),
      .ADR1 (\bridge/configuration/C1941 ),
      .ADR2 (\bridge/configuration/wb_err_addr [0]),
      .ADR3 (\bridge/configuration/wb_error_en ),
      .O (\syn179848/FROM )
    );
    X_BUF \syn179848/YUSED (
      .I (\syn179848/GROM ),
      .O (syn180995)
    );
    X_BUF \syn179848/XUSED (
      .I (\syn179848/FROM ),
      .O (syn179848)
    );
    defparam C17904.INIT = 16'h20E3;
    X_LUT4 C17904(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C723 ),
      .ADR1 (ERR_I),
      .ADR2 (ACK_I),
      .ADR3 (syn19555),
      .O (\N12311/GROM )
    );
    defparam C18818.INIT = 16'hBA00;
    X_LUT4 C18818(
      .ADR0 (syn19555),
      .ADR1 (ACK_I),
      .ADR2 (ERR_I),
      .ADR3 (syn179789),
      .O (\N12311/FROM )
    );
    X_BUF \N12311/YUSED (
      .I (\N12311/GROM ),
      .O (syn22790)
    );
    X_BUF \N12311/XUSED (
      .I (\N12311/FROM ),
      .O (N12311)
    );
    defparam C17760.INIT = 16'h9009;
    X_LUT4 C17760(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [4]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [4]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_next [3]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [3]),
      .O (\syn182394/GROM )
    );
    defparam C17763.INIT = 16'h7BDE;
    X_LUT4 C17763(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [4]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [4]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [3]),
      .O (\syn182394/FROM )
    );
    X_BUF \syn182394/YUSED (
      .I (\syn182394/GROM ),
      .O (syn182403)
    );
    X_BUF \syn182394/XUSED (
      .I (\syn182394/FROM ),
      .O (syn182394)
    );
    defparam C17744.INIT = 16'h9009;
    X_LUT4 C17744(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [2]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [2]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [1]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [1]),
      .O (\syn182432/GROM )
    );
    X_BUF \syn182432/YUSED (
      .I (\syn182432/GROM ),
      .O (syn182432)
    );
    defparam C19265.INIT = 16'hFA0A;
    X_LUT4 C19265(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_addr_out [16]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[16]/GROM )
    );
    defparam C19369.INIT = 16'hEEEE;
    X_LUT4 C19369(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[16]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<16>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[16]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [16])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<16>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[16]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [16])
    );
    defparam C19193.INIT = 16'hF0AA;
    X_LUT4 C19193(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pcit_if_addr_out [7]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[7]/GROM )
    );
    defparam C19336.INIT = 16'hFAFA;
    X_LUT4 C19336(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[7]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<7>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[7]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [7])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<7>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[7]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [7])
    );
    defparam C19185.INIT = 16'hCCA0;
    X_LUT4 C19185(
      .ADR0 (\CRT/pix_start_addr [15]),
      .ADR1 (\CRT/wbs_pal_data [15]),
      .ADR2 (ADR_O[2]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[31]/GROM )
    );
    defparam C19234.INIT = 16'h00A0;
    X_LUT4 C19234(
      .ADR0 (ADR_O[2]),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [31]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[31]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<31>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[31]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [15])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<31>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[31]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [31])
    );
    defparam C19177.INIT = 16'hE2C0;
    X_LUT4 C19177(
      .ADR0 (\CRT/pix_start_addr [7]),
      .ADR1 (ADR_O[10]),
      .ADR2 (\CRT/wbs_pal_data [7]),
      .ADR3 (ADR_O[2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[23]/GROM )
    );
    defparam C19226.INIT = 16'h0A00;
    X_LUT4 C19226(
      .ADR0 (\CRT/pix_start_addr [23]),
      .ADR1 (VCC),
      .ADR2 (ADR_O[10]),
      .ADR3 (ADR_O[2]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[23]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<23>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[23]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [7])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<23>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[23]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [23])
    );
    defparam C18617.INIT = 16'hECA0;
    X_LUT4 C18617(
      .ADR0 (\bridge/configuration/pci_err_addr [11]),
      .ADR1 (\bridge/configuration/pci_err_data [11]),
      .ADR2 (syn17107),
      .ADR3 (syn17109),
      .O (\syn180122/GROM )
    );
    defparam C18674.INIT = 16'hF888;
    X_LUT4 C18674(
      .ADR0 (syn17107),
      .ADR1 (\bridge/configuration/pci_err_addr [7]),
      .ADR2 (\bridge/configuration/pci_err_data [7]),
      .ADR3 (syn17109),
      .O (\syn180122/FROM )
    );
    X_BUF \syn180122/YUSED (
      .I (\syn180122/GROM ),
      .O (syn180284)
    );
    X_BUF \syn180122/XUSED (
      .I (\syn180122/FROM ),
      .O (syn180122)
    );
    defparam C18561.INIT = 16'hECA0;
    X_LUT4 C18561(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [14]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [14]),
      .ADR2 (syn16919),
      .ADR3 (syn16931),
      .O (\syn120384/GROM )
    );
    X_BUF \syn120384/YUSED (
      .I (\syn120384/GROM ),
      .O (syn120384)
    );
    defparam C18537.INIT = 16'hEC00;
    X_LUT4 C18537(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/configuration/C1953 ),
      .ADR2 (\bridge/configuration/wb_base_addr1 [16]),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [16]),
      .O (\syn178092/GROM )
    );
    defparam C19680.INIT = 16'hF8F0;
    X_LUT4 C19680(
      .ADR0 (\bridge/configuration/C2322 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [16]),
      .ADR2 (\bridge/configuration/C2368 ),
      .ADR3 (\bridge/configuration/wb_base_addr1 [16]),
      .O (\syn178092/FROM )
    );
    X_BUF \syn178092/YUSED (
      .I (\syn178092/GROM ),
      .O (syn21014)
    );
    X_BUF \syn178092/XUSED (
      .I (\syn178092/FROM ),
      .O (syn178092)
    );
    defparam C18529.INIT = 16'hE040;
    X_LUT4 C18529(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [16]),
      .ADR2 (syn19366),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [16]),
      .O (\syn120382/GROM )
    );
    defparam C18597.INIT = 16'hC480;
    X_LUT4 C18597(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .ADR1 (syn19366),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [12]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [12]),
      .O (\syn120382/FROM )
    );
    X_BUF \syn120382/YUSED (
      .I (\syn120382/GROM ),
      .O (syn180532)
    );
    X_BUF \syn120382/XUSED (
      .I (\syn120382/FROM ),
      .O (syn120382)
    );
    defparam C18377.INIT = 16'hF888;
    X_LUT4 C18377(
      .ADR0 (\bridge/configuration/wb_err_data [26]),
      .ADR1 (\bridge/configuration/C1935 ),
      .ADR2 (\bridge/conf_pci_ba0_out [14]),
      .ADR3 (\bridge/configuration/C2003 ),
      .O (\syn20770/GROM )
    );
    defparam C18644.INIT = 16'hA000;
    X_LUT4 C18644(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/configuration/wb_err_data [9]),
      .O (\syn20770/FROM )
    );
    X_BUF \syn20770/YUSED (
      .I (\syn20770/GROM ),
      .O (syn180994)
    );
    X_BUF \syn20770/XUSED (
      .I (\syn20770/FROM ),
      .O (syn20770)
    );
    defparam C17745.INIT = 16'h8241;
    X_LUT4 C17745(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [4]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_minus1 [3]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [3]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [4]),
      .O (\syn182423/GROM )
    );
    defparam C17748.INIT = 16'h9009;
    X_LUT4 C17748(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [4]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [4]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [3]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rgrey_addr [3]),
      .O (\syn182423/FROM )
    );
    X_BUF \syn182423/YUSED (
      .I (\syn182423/GROM ),
      .O (syn182431)
    );
    X_BUF \syn182423/XUSED (
      .I (\syn182423/FROM ),
      .O (syn182423)
    );
    defparam C19610.INIT = 16'hEAC0;
    X_LUT4 C19610(
      .ADR0 (\bridge/configuration/pci_base_addr0 [12]),
      .ADR1 (syn17067),
      .ADR2 (\bridge/conf_latency_tim_out [4]),
      .ADR3 (syn16930),
      .O (\syn178179/GROM )
    );
    defparam C19638.INIT = 16'hECA0;
    X_LUT4 C19638(
      .ADR0 (syn17067),
      .ADR1 (\bridge/configuration/pci_base_addr0 [14]),
      .ADR2 (\bridge/conf_latency_tim_out [6]),
      .ADR3 (syn16930),
      .O (\syn178179/FROM )
    );
    X_BUF \syn178179/YUSED (
      .I (\syn178179/GROM ),
      .O (syn178250)
    );
    X_BUF \syn178179/XUSED (
      .I (\syn178179/FROM ),
      .O (syn178179)
    );
    defparam C19530.INIT = 16'hEAEA;
    X_LUT4 C19530(
      .ADR0 (syn24326),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [3]),
      .ADR2 (syn17745),
      .ADR3 (VCC),
      .O (\syn24474/GROM )
    );
    defparam C19544.INIT = 16'hF8F8;
    X_LUT4 C19544(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [5]),
      .ADR1 (syn17745),
      .ADR2 (syn24326),
      .ADR3 (VCC),
      .O (\syn24474/FROM )
    );
    X_BUF \syn24474/YUSED (
      .I (\syn24474/GROM ),
      .O (syn24476)
    );
    X_BUF \syn24474/XUSED (
      .I (\syn24474/FROM ),
      .O (syn24474)
    );
    defparam C19274.INIT = 16'hCCF0;
    X_LUT4 C19274(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [25]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[25]/GROM )
    );
    defparam C19378.INIT = 16'hEEEE;
    X_LUT4 C19378(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[25]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<25>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[25]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [25])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<25>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[25]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [25])
    );
    defparam C19266.INIT = 16'hD8D8;
    X_LUT4 C19266(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [17]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[17]/GROM )
    );
    defparam C19370.INIT = 16'hEEEE;
    X_LUT4 C19370(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[17]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<17>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[17]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [17])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<17>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[17]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [17])
    );
    defparam C19194.INIT = 16'hD8D8;
    X_LUT4 C19194(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [8]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[8]/GROM )
    );
    defparam C19337.INIT = 16'hFFF0;
    X_LUT4 C19337(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[8]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<8>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[8]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [8])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<8>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[8]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [8])
    );
    defparam C19186.INIT = 16'hF5A0;
    X_LUT4 C19186(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pcit_if_addr_out [0]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .O (\bridge/pci_target_unit/pci_target_sm/S_291/cell0/GROM )
    );
    defparam C19303.INIT = 16'h1111;
    X_LUT4 C19303(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/in_reg_irdy_out ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/pci_target_sm/S_291/cell0/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/S_291/cell0/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/S_291/cell0/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [0])
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/S_291/cell0/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/S_291/cell0/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 )
    );
    defparam C19178.INIT = 16'hCAC0;
    X_LUT4 C19178(
      .ADR0 (ADR_O[2]),
      .ADR1 (\CRT/wbs_pal_data [8]),
      .ADR2 (ADR_O[10]),
      .ADR3 (\CRT/pix_start_addr [8]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[24]/GROM )
    );
    defparam C19227.INIT = 16'h00A0;
    X_LUT4 C19227(
      .ADR0 (ADR_O[2]),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [24]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[24]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<24>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[24]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [8])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<24>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[24]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [24])
    );
    defparam C18642.INIT = 16'hA000;
    X_LUT4 C18642(
      .ADR0 (\bridge/configuration/pci_err_data [9]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/configuration/C1967 ),
      .O (\syn16934/GROM )
    );
    defparam C18837.INIT = 16'h0C0C;
    X_LUT4 C18837(
      .ADR0 (VCC),
      .ADR1 (syn60111),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (VCC),
      .O (\syn16934/FROM )
    );
    X_BUF \syn16934/YUSED (
      .I (\syn16934/GROM ),
      .O (syn20772)
    );
    X_BUF \syn16934/XUSED (
      .I (\syn16934/FROM ),
      .O (syn16934)
    );
    defparam C18634.INIT = 16'hF888;
    X_LUT4 C18634(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [9]),
      .ADR1 (syn136384),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [9]),
      .ADR3 (syn136386),
      .O (\syn180098/GROM )
    );
    defparam C18680.INIT = 16'hEAC0;
    X_LUT4 C18680(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [6]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [6]),
      .ADR2 (syn136384),
      .ADR3 (syn136386),
      .O (\syn180098/FROM )
    );
    X_BUF \syn180098/YUSED (
      .I (\syn180098/GROM ),
      .O (syn180222)
    );
    X_BUF \syn180098/XUSED (
      .I (\syn180098/FROM ),
      .O (syn180098)
    );
    defparam C18618.INIT = 16'hEAC0;
    X_LUT4 C18618(
      .ADR0 (syn17110),
      .ADR1 (\bridge/configuration/wb_err_data [11]),
      .ADR2 (syn17111),
      .ADR3 (\bridge/configuration/wb_err_addr [11]),
      .O (\syn180121/GROM )
    );
    defparam C18675.INIT = 16'hEAC0;
    X_LUT4 C18675(
      .ADR0 (syn17110),
      .ADR1 (\bridge/configuration/wb_err_data [7]),
      .ADR2 (syn17111),
      .ADR3 (\bridge/configuration/wb_err_addr [7]),
      .O (\syn180121/FROM )
    );
    X_BUF \syn180121/YUSED (
      .I (\syn180121/GROM ),
      .O (syn180283)
    );
    X_BUF \syn180121/XUSED (
      .I (\syn180121/FROM ),
      .O (syn180121)
    );
    defparam C18490.INIT = 16'hC888;
    X_LUT4 C18490(
      .ADR0 (\bridge/configuration/C1953 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [19]),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/configuration/wb_base_addr1 [19]),
      .O (\syn21091/GROM )
    );
    defparam C18505.INIT = 16'hF800;
    X_LUT4 C18505(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/configuration/wb_base_addr1 [18]),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/configuration/wb_addr_mask1 [18]),
      .O (\syn21091/FROM )
    );
    X_BUF \syn21091/YUSED (
      .I (\syn21091/GROM ),
      .O (syn21130)
    );
    X_BUF \syn21091/XUSED (
      .I (\syn21091/FROM ),
      .O (syn21091)
    );
    defparam C18394.INIT = 16'hC888;
    X_LUT4 C18394(
      .ADR0 (\bridge/configuration/C1953 ),
      .ADR1 (\bridge/conf_wb_am1_out [13]),
      .ADR2 (\bridge/conf_wb_ba1_out [13]),
      .ADR3 (\bridge/configuration/C1955 ),
      .O (\syn60044/GROM )
    );
    defparam C19967.INIT = 16'hAF5F;
    X_LUT4 C19967(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [25]),
      .ADR1 (VCC),
      .ADR2 (\bridge/conf_wb_am1_out [13]),
      .ADR3 (\bridge/conf_wb_ba1_out [13]),
      .O (\syn60044/FROM )
    );
    X_BUF \syn60044/YUSED (
      .I (\syn60044/GROM ),
      .O (syn21365)
    );
    X_BUF \syn60044/XUSED (
      .I (\syn60044/FROM ),
      .O (syn60044)
    );
    defparam C19611.INIT = 16'hA000;
    X_LUT4 C19611(
      .ADR0 (syn16928),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/pci_base_addr1 [12]),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [12]),
      .O (\syn18468/GROM )
    );
    defparam C19639.INIT = 16'h8080;
    X_LUT4 C19639(
      .ADR0 (syn16928),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [14]),
      .ADR2 (\bridge/configuration/pci_base_addr1 [14]),
      .ADR3 (VCC),
      .O (\syn18468/FROM )
    );
    X_BUF \syn18468/YUSED (
      .I (\syn18468/GROM ),
      .O (syn18543)
    );
    X_BUF \syn18468/XUSED (
      .I (\syn18468/FROM ),
      .O (syn18468)
    );
    defparam C19515.INIT = 16'hEAC0;
    X_LUT4 C19515(
      .ADR0 (\bridge/configuration/pci_err_addr [2]),
      .ADR1 (\bridge/configuration/wb_err_data [2]),
      .ADR2 (\bridge/configuration/C2302 ),
      .ADR3 (\bridge/configuration/C2338 ),
      .O (\syn17071/GROM )
    );
    defparam C19606.INIT = 16'hAA00;
    X_LUT4 C19606(
      .ADR0 (syn16917),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C2338 ),
      .O (\syn17071/FROM )
    );
    X_BUF \syn17071/YUSED (
      .I (\syn17071/GROM ),
      .O (syn178460)
    );
    X_BUF \syn17071/XUSED (
      .I (\syn17071/FROM ),
      .O (syn17071)
    );
    defparam C19275.INIT = 16'hCFC0;
    X_LUT4 C19275(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [26]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[26]/GROM )
    );
    defparam C19379.INIT = 16'hFFAA;
    X_LUT4 C19379(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[26]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<26>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[26]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [26])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<26>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[26]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [26])
    );
    defparam C19267.INIT = 16'hB8B8;
    X_LUT4 C19267(
      .ADR0 (\bridge/pci_target_unit/pcit_if_addr_out [18]),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[18]/GROM )
    );
    defparam C19371.INIT = 16'hEEEE;
    X_LUT4 C19371(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[18]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<18>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[18]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [18])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<18>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[18]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [18])
    );
    defparam C19195.INIT = 16'hFC0C;
    X_LUT4 C19195(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [9]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_addr_out [9]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[9]/GROM )
    );
    defparam C19338.INIT = 16'hFFCC;
    X_LUT4 C19338(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [9]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[9]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<9>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[9]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [9])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<9>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[9]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [9])
    );
    defparam C19187.INIT = 16'hCACA;
    X_LUT4 C19187(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [1]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[1]/GROM )
    );
    defparam C19330.INIT = 16'hFCFC;
    X_LUT4 C19330(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[1]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<1>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[1]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [1])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<1>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[1]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [1])
    );
    defparam C19179.INIT = 16'hCCA0;
    X_LUT4 C19179(
      .ADR0 (\CRT/pix_start_addr [9]),
      .ADR1 (\CRT/wbs_pal_data [9]),
      .ADR2 (ADR_O[2]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[25]/GROM )
    );
    defparam C19228.INIT = 16'h00A0;
    X_LUT4 C19228(
      .ADR0 (ADR_O[2]),
      .ADR1 (VCC),
      .ADR2 (\CRT/pix_start_addr [25]),
      .ADR3 (ADR_O[10]),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[25]/FROM )
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<25>/YUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[25]/GROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [9])
    );
    X_BUF \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out<25>/XUSED (
      .I (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out[25]/FROM ),
      .O (\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [25])
    );
    defparam C18643.INIT = 16'h8080;
    X_LUT4 C18643(
      .ADR0 (\bridge/configuration/wb_err_addr [9]),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1937 ),
      .ADR3 (VCC),
      .O (\syn17102/GROM )
    );
    defparam C18732.INIT = 16'h2200;
    X_LUT4 C18732(
      .ADR0 (\bridge/configuration/C2268 ),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (VCC),
      .ADR3 (syn60111),
      .O (\syn17102/FROM )
    );
    X_BUF \syn17102/YUSED (
      .I (\syn17102/GROM ),
      .O (syn20771)
    );
    X_BUF \syn17102/XUSED (
      .I (\syn17102/FROM ),
      .O (syn17102)
    );
    defparam C18627.INIT = 16'h8800;
    X_LUT4 C18627(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/configuration/pci_err_addr [10]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\syn20773/GROM )
    );
    defparam C18641.INIT = 16'h8800;
    X_LUT4 C18641(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (\bridge/configuration/pci_err_addr [9]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\syn20773/FROM )
    );
    X_BUF \syn20773/YUSED (
      .I (\syn20773/GROM ),
      .O (syn20803)
    );
    X_BUF \syn20773/XUSED (
      .I (\syn20773/FROM ),
      .O (syn20773)
    );
    defparam C18547.INIT = 16'hECA0;
    X_LUT4 C18547(
      .ADR0 (\bridge/configuration/pci_err_data [15]),
      .ADR1 (\bridge/configuration/C1971 ),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (\bridge/configuration/pci_err_addr [15]),
      .O (\syn180420/GROM )
    );
    defparam C18564.INIT = 16'hEAC0;
    X_LUT4 C18564(
      .ADR0 (\bridge/configuration/pci_err_data [14]),
      .ADR1 (\bridge/configuration/pci_err_addr [14]),
      .ADR2 (\bridge/configuration/C1971 ),
      .ADR3 (\bridge/configuration/C1967 ),
      .O (\syn180420/FROM )
    );
    X_BUF \syn180420/YUSED (
      .I (\syn180420/GROM ),
      .O (syn180470)
    );
    X_BUF \syn180420/XUSED (
      .I (\syn180420/FROM ),
      .O (syn180420)
    );
    defparam C18299.INIT = 16'hF888;
    X_LUT4 C18299(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [30]),
      .ADR2 (syn17051),
      .ADR3 (syn60110),
      .O (\syn181037/GROM )
    );
    defparam C18355.INIT = 16'hEAC0;
    X_LUT4 C18355(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (syn17054),
      .ADR2 (syn60110),
      .ADR3 (\bridge/configuration/wb_tran_addr1 [27]),
      .O (\syn181037/FROM )
    );
    X_BUF \syn181037/YUSED (
      .I (\syn181037/GROM ),
      .O (syn181193)
    );
    X_BUF \syn181037/XUSED (
      .I (\syn181037/FROM ),
      .O (syn181037)
    );
    defparam C17691.INIT = 16'h6FF6;
    X_LUT4 C17691(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [3]),
      .O (\syn182526/GROM )
    );
    X_BUF \syn182526/YUSED (
      .I (\syn182526/GROM ),
      .O (syn182526)
    );
    defparam C19620.INIT = 16'hF888;
    X_LUT4 C19620(
      .ADR0 (\bridge/configuration/C2318 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [12]),
      .ADR2 (\bridge/configuration/wb_err_data [12]),
      .ADR3 (\bridge/configuration/C2302 ),
      .O (\syn178201/GROM )
    );
    defparam C19634.INIT = 16'hF888;
    X_LUT4 C19634(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [13]),
      .ADR1 (\bridge/configuration/C2318 ),
      .ADR2 (\bridge/configuration/wb_err_data [13]),
      .ADR3 (\bridge/configuration/C2302 ),
      .O (\syn178201/FROM )
    );
    X_BUF \syn178201/YUSED (
      .I (\syn178201/GROM ),
      .O (syn178237)
    );
    X_BUF \syn178201/XUSED (
      .I (\syn178201/FROM ),
      .O (syn178201)
    );
    defparam C19276.INIT = 16'hCCAA;
    X_LUT4 C19276(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [27]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[28]/GROM )
    );
    defparam C19277.INIT = 16'hAAF0;
    X_LUT4 C19277(
      .ADR0 (\bridge/pci_target_unit/pcit_if_addr_out [28]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[28]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<28>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[28]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [27])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<28>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[28]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [28])
    );
    defparam C19268.INIT = 16'hFC30;
    X_LUT4 C19268(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .ADR3 (\bridge/pci_target_unit/pcit_if_addr_out [19]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[20]/GROM )
    );
    defparam C19269.INIT = 16'hAAF0;
    X_LUT4 C19269(
      .ADR0 (\bridge/pci_target_unit/pcit_if_addr_out [20]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[20]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<20>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[20]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [19])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<20>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[20]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [20])
    );
    defparam C19196.INIT = 16'hD8D8;
    X_LUT4 C19196(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [10]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [10]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[10]/GROM )
    );
    defparam C19339.INIT = 16'hFFCC;
    X_LUT4 C19339(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [10]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[10]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<10>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[10]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [10])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<10>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[10]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [10])
    );
    defparam C19188.INIT = 16'hDD88;
    X_LUT4 C19188(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [2]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[2]/GROM )
    );
    defparam C19331.INIT = 16'hEEEE;
    X_LUT4 C19331(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[2]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<2>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[2]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [2])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<2>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[2]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [2])
    );
    defparam C18724.INIT = 16'hF888;
    X_LUT4 C18724(
      .ADR0 (\bridge/configuration/pci_err_data [3]),
      .ADR1 (syn16985),
      .ADR2 (\bridge/configuration/wb_err_addr [3]),
      .ADR3 (syn17014),
      .O (\syn178436/GROM )
    );
    defparam C19525.INIT = 16'hECA0;
    X_LUT4 C19525(
      .ADR0 (syn17081),
      .ADR1 (syn17077),
      .ADR2 (\bridge/conf_cache_line_size_out [3]),
      .ADR3 (\bridge/configuration/pci_err_data [3]),
      .O (\syn178436/FROM )
    );
    X_BUF \syn178436/YUSED (
      .I (\syn178436/GROM ),
      .O (syn179988)
    );
    X_BUF \syn178436/XUSED (
      .I (\syn178436/FROM ),
      .O (syn178436)
    );
    defparam C18708.INIT = 16'h8888;
    X_LUT4 C18708(
      .ADR0 (\bridge/configuration/C1971 ),
      .ADR1 (syn16916),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn179850/GROM )
    );
    defparam C18797.INIT = 16'hF888;
    X_LUT4 C18797(
      .ADR0 (\bridge/configuration/pci_err_addr [0]),
      .ADR1 (\bridge/configuration/C1971 ),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (\bridge/configuration/pci_err_data [0]),
      .O (\syn179850/FROM )
    );
    X_BUF \syn179850/YUSED (
      .I (\syn179850/GROM ),
      .O (syn17107)
    );
    X_BUF \syn179850/XUSED (
      .I (\syn179850/FROM ),
      .O (syn179850)
    );
    defparam C18660.INIT = 16'h8000;
    X_LUT4 C18660(
      .ADR0 (\bridge/conf_serr_enable_out ),
      .ADR1 (syn60038),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn17099),
      .O (\syn21507/GROM )
    );
    defparam C18327.INIT = 16'h8000;
    X_LUT4 C18327(
      .ADR0 (\bridge/conf_pci_ba1_out [16]),
      .ADR1 (\bridge/conf_pci_am1_out [16]),
      .ADR2 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR3 (syn16927),
      .O (\syn21507/FROM )
    );
    X_BUF \syn21507/YUSED (
      .I (\syn21507/GROM ),
      .O (syn20737)
    );
    X_BUF \syn21507/XUSED (
      .I (\syn21507/FROM ),
      .O (syn21507)
    );
    defparam C17908.INIT = 16'h0055;
    X_LUT4 C17908(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/c_state [0]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/c_state [1]),
      .O (\bridge/pci_target_unit/wishbone_master/C983/GROM )
    );
    defparam C19257.INIT = 16'h0011;
    X_LUT4 C19257(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/c_state [0]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/c_state [2]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/c_state [1]),
      .O (\bridge/pci_target_unit/wishbone_master/C983/FROM )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/C983/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/C983/GROM ),
      .O (syn19580)
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/C983/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/C983/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C983 )
    );
    defparam C17676.INIT = 16'h8241;
    X_LUT4 C17676(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [3]),
      .O (\syn182535/GROM )
    );
    defparam C17688.INIT = 16'h8241;
    X_LUT4 C17688(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_next [4]),
      .O (\syn182535/FROM )
    );
    X_BUF \syn182535/YUSED (
      .I (\syn182535/GROM ),
      .O (syn182564)
    );
    X_BUF \syn182535/XUSED (
      .I (\syn182535/FROM ),
      .O (syn182535)
    );
    defparam C17668.INIT = 16'h8421;
    X_LUT4 C17668(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [4]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_minus2 [4]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [3]),
      .O (\syn182555/GROM )
    );
    defparam C17673.INIT = 16'h8421;
    X_LUT4 C17673(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [3]),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [4]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [3]),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/rgrey_addr [4]),
      .O (\syn182555/FROM )
    );
    X_BUF \syn182555/YUSED (
      .I (\syn182555/GROM ),
      .O (syn182576)
    );
    X_BUF \syn182555/XUSED (
      .I (\syn182555/FROM ),
      .O (syn182555)
    );
    defparam C19437.INIT = 16'hF000;
    X_LUT4 C19437(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [2])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .O (\syn18965/GROM )
    );
    defparam C19440.INIT = 16'hF000;
    X_LUT4 C19440(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/raddr_plus_one [3])
      ,
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/rallow ),
      .O (\syn18965/FROM )
    );
    X_BUF \syn18965/YUSED (
      .I (\syn18965/GROM ),
      .O (syn18972)
    );
    X_BUF \syn18965/XUSED (
      .I (\syn18965/FROM ),
      .O (syn18965)
    );
    defparam C19373.INIT = 16'hFCFC;
    X_LUT4 C19373(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[22]/GROM )
    );
    defparam C19375.INIT = 16'hFFCC;
    X_LUT4 C19375(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[22]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<22>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[22]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [20])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<22>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[22]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [22])
    );
    defparam C17933.INIT = 16'hCC80;
    X_LUT4 C17933(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C983 ),
      .ADR1 (\bridge/pci_target_unit/fifos_pciw_control_out [0]),
      .ADR2 (syn17011),
      .ADR3 (syn179021),
      .O (\bridge/pci_target_unit/fifos/out_count_en/GROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/out_count_en/YUSED (
      .I (\bridge/pci_target_unit/fifos/out_count_en/GROM ),
      .O (\bridge/pci_target_unit/fifos/out_count_en )
    );
    defparam C19197.INIT = 16'hFC0C;
    X_LUT4 C19197(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [11]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_addr_out [11]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[12]/GROM )
    );
    defparam C19198.INIT = 16'hFC0C;
    X_LUT4 C19198(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_addr_out [12]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[12]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<12>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[12]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [11])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<12>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[12]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [12])
    );
    defparam C19189.INIT = 16'hEE44;
    X_LUT4 C19189(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pcit_if_addr_out [3]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[3]/GROM )
    );
    defparam C19332.INIT = 16'hFFCC;
    X_LUT4 C19332(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[3]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<3>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[3]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [3])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<3>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[3]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [3])
    );
    defparam C18813.INIT = 16'h0080;
    X_LUT4 C18813(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1925 ),
      .ADR3 (\bridge/in_reg_cbe_out [0]),
      .O (\bridge/configuration/C292/N3/GROM )
    );
    defparam C18822.INIT = 16'h4000;
    X_LUT4 C18822(
      .ADR0 (\bridge/in_reg_cbe_out [0]),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1973 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C292/N3/FROM )
    );
    X_BUF \bridge/configuration/C292/N3/YUSED (
      .I (\bridge/configuration/C292/N3/GROM ),
      .O (\bridge/configuration/C302/N19 )
    );
    X_BUF \bridge/configuration/C292/N3/XUSED (
      .I (\bridge/configuration/C292/N3/FROM ),
      .O (\bridge/configuration/C292/N3 )
    );
    defparam C18717.INIT = 16'hECA0;
    X_LUT4 C18717(
      .ADR0 (syn136386),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [3]),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [3]),
      .ADR3 (syn136384),
      .O (\syn179878/GROM )
    );
    defparam C18767.INIT = 16'hF888;
    X_LUT4 C18767(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_data_out [0]),
      .ADR1 (syn136386),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [0]),
      .ADR3 (syn136384),
      .O (\syn179878/FROM )
    );
    X_BUF \syn179878/YUSED (
      .I (\syn179878/GROM ),
      .O (syn180003)
    );
    X_BUF \syn179878/XUSED (
      .I (\syn179878/FROM ),
      .O (syn179878)
    );
    defparam C18653.INIT = 16'h8000;
    X_LUT4 C18653(
      .ADR0 (syn60038),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn17014),
      .ADR3 (\bridge/configuration/wb_err_addr [8]),
      .O (\syn20740/GROM )
    );
    defparam C18654.INIT = 16'h8000;
    X_LUT4 C18654(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (syn17015),
      .ADR2 (syn60038),
      .ADR3 (\bridge/configuration/wb_err_data [8]),
      .O (\syn20740/FROM )
    );
    X_BUF \syn20740/YUSED (
      .I (\syn20740/GROM ),
      .O (syn20741)
    );
    X_BUF \syn20740/XUSED (
      .I (\syn20740/FROM ),
      .O (syn20740)
    );
    defparam C18565.INIT = 16'hEAC0;
    X_LUT4 C18565(
      .ADR0 (\bridge/configuration/C1937 ),
      .ADR1 (\bridge/configuration/C1935 ),
      .ADR2 (\bridge/configuration/wb_err_data [14]),
      .ADR3 (\bridge/configuration/wb_err_addr [14]),
      .O (\syn179950/GROM )
    );
    defparam C18744.INIT = 16'hECA0;
    X_LUT4 C18744(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (\bridge/configuration/C1937 ),
      .ADR2 (\bridge/configuration/wb_err_data [2]),
      .ADR3 (\bridge/configuration/wb_err_addr [2]),
      .O (\syn179950/FROM )
    );
    X_BUF \syn179950/YUSED (
      .I (\syn179950/GROM ),
      .O (syn180419)
    );
    X_BUF \syn179950/XUSED (
      .I (\syn179950/FROM ),
      .O (syn179950)
    );
    defparam C18549.INIT = 16'hEAC0;
    X_LUT4 C18549(
      .ADR0 (\bridge/configuration/C2003 ),
      .ADR1 (\bridge/configuration/C1929 ),
      .ADR2 (\bridge/configuration/config_addr[15] ),
      .ADR3 (\bridge/configuration/pci_base_addr0 [15]),
      .O (\syn20769/GROM )
    );
    defparam C18637.INIT = 16'hC000;
    X_LUT4 C18637(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/C1929 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/configuration/config_addr[9] ),
      .O (\syn20769/FROM )
    );
    X_BUF \syn20769/YUSED (
      .I (\syn20769/GROM ),
      .O (syn180468)
    );
    X_BUF \syn20769/XUSED (
      .I (\syn20769/FROM ),
      .O (syn20769)
    );
    defparam C18485.INIT = 16'hECA0;
    X_LUT4 C18485(
      .ADR0 (\bridge/configuration/pci_err_data [19]),
      .ADR1 (\bridge/configuration/pci_err_addr [19]),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (\bridge/configuration/C1971 ),
      .O (\syn180611/GROM )
    );
    defparam C18500.INIT = 16'hF888;
    X_LUT4 C18500(
      .ADR0 (\bridge/configuration/pci_err_addr [18]),
      .ADR1 (\bridge/configuration/C1971 ),
      .ADR2 (\bridge/configuration/C1967 ),
      .ADR3 (\bridge/configuration/pci_err_data [18]),
      .O (\syn180611/FROM )
    );
    X_BUF \syn180611/YUSED (
      .I (\syn180611/GROM ),
      .O (syn180661)
    );
    X_BUF \syn180611/XUSED (
      .I (\syn180611/FROM ),
      .O (syn180611)
    );
    defparam C19630.INIT = 16'hF888;
    X_LUT4 C19630(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [13]),
      .ADR1 (\bridge/configuration/C2354 ),
      .ADR2 (\bridge/configuration/C2356 ),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [13]),
      .O (\syn177820/GROM )
    );
    defparam C19783.INIT = 16'hF888;
    X_LUT4 C19783(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [24]),
      .ADR1 (\bridge/configuration/C2354 ),
      .ADR2 (\bridge/conf_pci_am1_out [12]),
      .ADR3 (\bridge/configuration/C2356 ),
      .O (\syn177820/FROM )
    );
    X_BUF \syn177820/YUSED (
      .I (\syn177820/GROM ),
      .O (syn178207)
    );
    X_BUF \syn177820/XUSED (
      .I (\syn177820/FROM ),
      .O (syn177820)
    );
    defparam C19454.INIT = 16'hFFEE;
    X_LUT4 C19454(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .ADR1 (N12359),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/load_force/GROM )
    );
    defparam C19473.INIT = 16'hEECC;
    X_LUT4 C19473(
      .ADR0 (N12359),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 ),
      .ADR2 (VCC),
      .ADR3 (syn17023),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/load_force/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/load_force/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/load_force/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/frame_load_slow )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/load_force/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/load_force/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/load_force )
    );
    defparam C19446.INIT = 16'hFFDD;
    X_LUT4 C19446(
      .ADR0 (syn16935),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/empty ),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/stretched_empty ),
      .O (\syn18944/GROM )
    );
    X_BUF \syn18944/YUSED (
      .I (\syn18944/GROM ),
      .O (syn18944)
    );
    defparam C19278.INIT = 16'hAAF0;
    X_LUT4 C19278(
      .ADR0 (\bridge/pci_target_unit/pcit_if_addr_out [29]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[30]/GROM )
    );
    defparam C19279.INIT = 16'hCCF0;
    X_LUT4 C19279(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_if_addr_out [30]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[30]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<30>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[30]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [29])
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out<30>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out[30]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [30])
    );
    defparam C18902.INIT = 16'h4000;
    X_LUT4 C18902(
      .ADR0 (\bridge/in_reg_cbe_out [0]),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/pci_target_unit/pci_target_if/n_1298/GROM )
    );
    defparam C19074.INIT = 16'hA000;
    X_LUT4 C19074(
      .ADR0 (\bridge/in_reg_cbe_out [2]),
      .ADR1 (VCC),
      .ADR2 (\bridge/in_reg_cbe_out [1]),
      .ADR3 (\bridge/in_reg_cbe_out [0]),
      .O (\bridge/pci_target_unit/pci_target_if/n_1298/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_if/n_1298/YUSED (
      .I (\bridge/pci_target_unit/pci_target_if/n_1298/GROM ),
      .O (\bridge/configuration/C299/N99 )
    );
    X_BUF \bridge/pci_target_unit/pci_target_if/n_1298/XUSED (
      .I (\bridge/pci_target_unit/pci_target_if/n_1298/FROM ),
      .O (\bridge/pci_target_unit/pci_target_if/n_1298 )
    );
    defparam C18830.INIT = 16'h0400;
    X_LUT4 C18830(
      .ADR0 (\bridge/pciu_conf_offset_out [3]),
      .ADR1 (\bridge/pciu_conf_offset_out [6]),
      .ADR2 (\bridge/in_reg_cbe_out [1]),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\bridge/configuration/C346/N5/GROM )
    );
    defparam C18857.INIT = 16'h4040;
    X_LUT4 C18857(
      .ADR0 (\bridge/in_reg_cbe_out [1]),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1941 ),
      .ADR3 (VCC),
      .O (\bridge/configuration/C346/N5/FROM )
    );
    X_BUF \bridge/configuration/C346/N5/YUSED (
      .I (\bridge/configuration/C346/N5/GROM ),
      .O (syn179775)
    );
    X_BUF \bridge/configuration/C346/N5/XUSED (
      .I (\bridge/configuration/C346/N5/FROM ),
      .O (\bridge/configuration/C346/N5 )
    );
    defparam C18806.INIT = 16'h2000;
    X_LUT4 C18806(
      .ADR0 (\bridge/configuration/C2268 ),
      .ADR1 (\bridge/in_reg_cbe_out [1]),
      .ADR2 (syn16934),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C284/N39/GROM )
    );
    defparam C18807.INIT = 16'h2000;
    X_LUT4 C18807(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/in_reg_cbe_out [0]),
      .ADR2 (\bridge/configuration/C2268 ),
      .ADR3 (syn16934),
      .O (\bridge/configuration/C284/N39/FROM )
    );
    X_BUF \bridge/configuration/C284/N39/YUSED (
      .I (\bridge/configuration/C284/N39/GROM ),
      .O (\bridge/configuration/C283/N39 )
    );
    X_BUF \bridge/configuration/C284/N39/XUSED (
      .I (\bridge/configuration/C284/N39/FROM ),
      .O (\bridge/configuration/C284/N39 )
    );
    defparam C18742.INIT = 16'hECA0;
    X_LUT4 C18742(
      .ADR0 (\bridge/configuration/C1967 ),
      .ADR1 (\bridge/configuration/wb_img_ctrl1[2] ),
      .ADR2 (\bridge/configuration/pci_err_data [2]),
      .ADR3 (\bridge/configuration/C1959 ),
      .O (\syn179912/GROM )
    );
    defparam C18756.INIT = 16'hECA0;
    X_LUT4 C18756(
      .ADR0 (\bridge/configuration/C1937 ),
      .ADR1 (\bridge/configuration/C1959 ),
      .ADR2 (\bridge/configuration/wb_err_addr [1]),
      .ADR3 (\bridge/conf_wb_img_ctrl1_out [1]),
      .O (\syn179912/FROM )
    );
    X_BUF \syn179912/YUSED (
      .I (\syn179912/GROM ),
      .O (syn179951)
    );
    X_BUF \syn179912/XUSED (
      .I (\syn179912/FROM ),
      .O (syn179912)
    );
    defparam C18590.INIT = 16'hE0C0;
    X_LUT4 C18590(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/configuration/C1953 ),
      .ADR2 (\bridge/configuration/wb_addr_mask1 [13]),
      .ADR3 (\bridge/configuration/wb_base_addr1 [13]),
      .O (\syn178200/GROM )
    );
    defparam C19635.INIT = 16'hF8F0;
    X_LUT4 C19635(
      .ADR0 (\bridge/configuration/wb_addr_mask1 [13]),
      .ADR1 (\bridge/configuration/C2322 ),
      .ADR2 (\bridge/configuration/C2368 ),
      .ADR3 (\bridge/configuration/wb_base_addr1 [13]),
      .O (\syn178200/FROM )
    );
    X_BUF \syn178200/YUSED (
      .I (\syn178200/GROM ),
      .O (syn20893)
    );
    X_BUF \syn178200/XUSED (
      .I (\syn178200/FROM ),
      .O (syn178200)
    );
    defparam C18398.INIT = 16'hECA0;
    X_LUT4 C18398(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [24]),
      .ADR1 (syn16919),
      .ADR2 (syn16931),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [24]),
      .O (\syn120386/GROM )
    );
    defparam C18544.INIT = 16'hECA0;
    X_LUT4 C18544(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [15]),
      .ADR1 (syn16919),
      .ADR2 (syn16931),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [15]),
      .O (\syn120386/FROM )
    );
    X_BUF \syn120386/YUSED (
      .I (\syn120386/GROM ),
      .O (syn120394)
    );
    X_BUF \syn120386/XUSED (
      .I (\syn120386/FROM ),
      .O (syn120386)
    );
    defparam C17950.INIT = 16'h8241;
    X_LUT4 C17950(
      .ADR0 (\bridge/pci_target_unit/del_sync_bc_out [0]),
      .ADR1 (\bridge/pci_target_unit/del_sync_bc_out [3]),
      .ADR2 (\bridge/in_reg_cbe_out [3]),
      .ADR3 (\bridge/in_reg_cbe_out [0]),
      .O (\bridge/pci_target_unit/pci_target_if/n_1335/GROM )
    );
    defparam C19072.INIT = 16'hB030;
    X_LUT4 C19072(
      .ADR0 (\bridge/in_reg_cbe_out [2]),
      .ADR1 (\bridge/in_reg_cbe_out [1]),
      .ADR2 (\bridge/in_reg_cbe_out [0]),
      .ADR3 (\bridge/in_reg_cbe_out [3]),
      .O (\bridge/pci_target_unit/pci_target_if/n_1335/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_if/n_1335/YUSED (
      .I (\bridge/pci_target_unit/pci_target_if/n_1335/GROM ),
      .O (syn182005)
    );
    X_BUF \bridge/pci_target_unit/pci_target_if/n_1335/XUSED (
      .I (\bridge/pci_target_unit/pci_target_if/n_1335/FROM ),
      .O (\bridge/pci_target_unit/pci_target_if/n_1335 )
    );
    defparam C19535.INIT = 16'h8080;
    X_LUT4 C19535(
      .ADR0 (syn16917),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (\bridge/configuration/wb_err_data [4]),
      .ADR3 (VCC),
      .O (\syn18655/GROM )
    );
    defparam C19558.INIT = 16'h8800;
    X_LUT4 C19558(
      .ADR0 (syn16917),
      .ADR1 (\bridge/configuration/wb_err_data [7]),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C2302 ),
      .O (\syn18655/FROM )
    );
    X_BUF \syn18655/YUSED (
      .I (\syn18655/GROM ),
      .O (syn18713)
    );
    X_BUF \syn18655/XUSED (
      .I (\syn18655/FROM ),
      .O (syn18655)
    );
    defparam C19199.INIT = 16'hF3C0;
    X_LUT4 C19199(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR2 (\bridge/pci_target_unit/pcit_if_addr_out [13]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[13]/GROM )
    );
    defparam C19342.INIT = 16'hFFCC;
    X_LUT4 C19342(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[13]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<13>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[13]/GROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [13])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<13>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[13]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [13])
    );
    defparam C18727.INIT = 16'hECA0;
    X_LUT4 C18727(
      .ADR0 (\bridge/configuration/wb_err_data [3]),
      .ADR1 (\bridge/configuration/config_addr[3] ),
      .ADR2 (syn17015),
      .ADR3 (syn17016),
      .O (\syn178433/GROM )
    );
    defparam C19523.INIT = 16'hECA0;
    X_LUT4 C19523(
      .ADR0 (\bridge/configuration/wb_err_addr [3]),
      .ADR1 (\bridge/configuration/config_addr[3] ),
      .ADR2 (syn17078),
      .ADR3 (syn17079),
      .O (\syn178433/FROM )
    );
    X_BUF \syn178433/YUSED (
      .I (\syn178433/GROM ),
      .O (syn179987)
    );
    X_BUF \syn178433/XUSED (
      .I (\syn178433/FROM ),
      .O (syn178433)
    );
    defparam C18647.INIT = 16'hECA0;
    X_LUT4 C18647(
      .ADR0 (syn20493),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_data_out [9]),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [9]),
      .O (\syn180107/GROM )
    );
    defparam C18671.INIT = 16'hEAC0;
    X_LUT4 C18671(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [7]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_data_out [7]),
      .ADR2 (syn20493),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .O (\syn180107/FROM )
    );
    X_BUF \syn180107/YUSED (
      .I (\syn180107/GROM ),
      .O (syn180219)
    );
    X_BUF \syn180107/XUSED (
      .I (\syn180107/FROM ),
      .O (syn180107)
    );
    defparam C18487.INIT = 16'hEAC0;
    X_LUT4 C18487(
      .ADR0 (\bridge/configuration/config_addr[19] ),
      .ADR1 (\bridge/configuration/C2003 ),
      .ADR2 (\bridge/configuration/pci_base_addr0 [19]),
      .ADR3 (\bridge/configuration/C1929 ),
      .O (\syn180609/GROM )
    );
    defparam C18502.INIT = 16'hF888;
    X_LUT4 C18502(
      .ADR0 (\bridge/configuration/pci_base_addr0 [18]),
      .ADR1 (\bridge/configuration/C2003 ),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/configuration/config_addr[18] ),
      .O (\syn180609/FROM )
    );
    X_BUF \syn180609/YUSED (
      .I (\syn180609/GROM ),
      .O (syn180659)
    );
    X_BUF \syn180609/XUSED (
      .I (\syn180609/FROM ),
      .O (syn180609)
    );
    defparam C17951.INIT = 16'h8421;
    X_LUT4 C17951(
      .ADR0 (\bridge/pci_target_unit/del_sync_bc_out [2]),
      .ADR1 (\bridge/in_reg_cbe_out [1]),
      .ADR2 (\bridge/in_reg_cbe_out [2]),
      .ADR3 (\bridge/pci_target_unit/del_sync_bc_out [1]),
      .O (\syn17031/GROM )
    );
    defparam C19319.INIT = 16'h3300;
    X_LUT4 C19319(
      .ADR0 (VCC),
      .ADR1 (\bridge/in_reg_cbe_out [2]),
      .ADR2 (VCC),
      .ADR3 (\bridge/in_reg_cbe_out [1]),
      .O (\syn17031/FROM )
    );
    X_BUF \syn17031/YUSED (
      .I (\syn17031/GROM ),
      .O (syn182004)
    );
    X_BUF \syn17031/XUSED (
      .I (\syn17031/FROM ),
      .O (syn17031)
    );
    defparam C17943.INIT = 16'h9009;
    X_LUT4 C17943(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [5]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [4]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[5]/GROM )
    );
    defparam C19334.INIT = 16'hFFAA;
    X_LUT4 C19334(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[5]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<5>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[5]/GROM ),
      .O (syn182001)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<5>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[5]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [5])
    );
    defparam C17919.INIT = 16'h20A0;
    X_LUT4 C17919(
      .ADR0 (\bridge/in_reg_frame_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/bckp_trdy_reg ),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/same_read_reg ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/trdy_asserted_reg ),
      .O (\syn17023/GROM )
    );
    defparam C19475.INIT = 16'h00C0;
    X_LUT4 C19475(
      .ADR0 (VCC),
      .ADR1 (\bridge/in_reg_irdy_out ),
      .ADR2 (\bridge/in_reg_frame_out ),
      .ADR3 (N_GNT),
      .O (\syn17023/FROM )
    );
    X_BUF \syn17023/YUSED (
      .I (\syn17023/GROM ),
      .O (syn182052)
    );
    X_BUF \syn17023/XUSED (
      .I (\syn17023/FROM ),
      .O (syn17023)
    );
    defparam C17783.INIT = 16'hA0A0;
    X_LUT4 C17783(
      .ADR0 (\bridge/pci_target_unit/del_sync/comp_rty_exp_clr ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg/GROM )
    );
    defparam C17784.INIT = 16'h33FF;
    X_LUT4 C17784(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/comp_rty_exp_clr ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg ),
      .O (N12602)
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_rty_exp_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/del_sync/comp_rty_exp_reg/YUSED (
      .I (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg/GROM ),
      .O (N12539)
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_rty_exp_reg_reg (
      .I (N12602),
      .CLK (CLK_BUFGPed),
      .CE (N12539),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_rty_exp_reg/FFX/ASYNC_FF_GSR_OR_145 (
      .I0 (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_rty_exp_reg/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19800.INIT = 16'hFEFA;
    X_LUT4 C19800(
      .ADR0 (syn24559),
      .ADR1 (syn17056),
      .ADR2 (syn18066),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn17895/GROM )
    );
    defparam C19867.INIT = 16'h8080;
    X_LUT4 C19867(
      .ADR0 (\bridge/conf_pci_ba1_out [17]),
      .ADR1 (\bridge/conf_pci_am1_out [17]),
      .ADR2 (\bridge/configuration/C2360 ),
      .ADR3 (VCC),
      .O (\syn17895/FROM )
    );
    X_BUF \syn17895/YUSED (
      .I (\syn17895/GROM ),
      .O (syn177780)
    );
    X_BUF \syn17895/XUSED (
      .I (\syn17895/FROM ),
      .O (syn17895)
    );
    defparam C19624.INIT = 16'hEAC0;
    X_LUT4 C19624(
      .ADR0 (\bridge/conf_latency_tim_out [5]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [13]),
      .ADR2 (syn17745),
      .ADR3 (syn17067),
      .O (\syn178106/GROM )
    );
    defparam C19667.INIT = 16'hEAC0;
    X_LUT4 C19667(
      .ADR0 (syn16930),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [16]),
      .ADR2 (syn17745),
      .ADR3 (\bridge/configuration/pci_base_addr0 [16]),
      .O (\syn178106/FROM )
    );
    X_BUF \syn178106/YUSED (
      .I (\syn178106/GROM ),
      .O (syn178214)
    );
    X_BUF \syn178106/XUSED (
      .I (\syn178106/FROM ),
      .O (syn178106)
    );
    defparam C19536.INIT = 16'hF888;
    X_LUT4 C19536(
      .ADR0 (\bridge/configuration/config_addr[4] ),
      .ADR1 (syn17076),
      .ADR2 (syn17073),
      .ADR3 (\bridge/configuration/wb_err_addr [4]),
      .O (\syn178356/GROM )
    );
    defparam C19559.INIT = 16'hEAC0;
    X_LUT4 C19559(
      .ADR0 (\bridge/configuration/wb_err_addr [7]),
      .ADR1 (syn17076),
      .ADR2 (\bridge/configuration/config_addr[7] ),
      .ADR3 (syn17073),
      .O (\syn178356/FROM )
    );
    X_BUF \syn178356/YUSED (
      .I (\syn178356/GROM ),
      .O (syn178409)
    );
    X_BUF \syn178356/XUSED (
      .I (\syn178356/FROM ),
      .O (syn178356)
    );
    defparam C19456.INIT = 16'h0008;
    X_LUT4 C19456(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .ADR1 (syn17010),
      .ADR2 (N_GNT),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/GROM )
    );
    defparam C18219.INIT = 16'h5D55;
    X_LUT4 C18219(
      .ADR0 (syn18858),
      .ADR1 (syn17010),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N40 )
    );
    X_INV \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<0>/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/GROM ),
      .O (syn18939)
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state_reg<0> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N40 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_sm/change_state ),
      .SET 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/FFX/ASYNC_FF_GSR_OR )
      ,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_sm/cur_state<0>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state[0]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19368.INIT = 16'h1111;
    X_LUT4 C19368(
      .ADR0 (N12360),
      .ADR1 (syn177324),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow/GROM )
    );
    defparam C19450.INIT = 16'h0101;
    X_LUT4 C19450(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_full_out ),
      .ADR1 (syn177324),
      .ADR2 (N12360),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow/GROM ),
      .O (\bridge/wishbone_slave_unit/wbs_sm_wbw_control_out [0])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow/FROM ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow )
    );
    defparam C18904.INIT = 16'h1111;
    X_LUT4 C18904(
      .ADR0 (\bridge/pciu_conf_offset_out [3]),
      .ADR1 (\bridge/pciu_conf_offset_out [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn17005/GROM )
    );
    X_BUF \syn17005/YUSED (
      .I (\syn17005/GROM ),
      .O (syn17005)
    );
    defparam C18832.INIT = 16'h3030;
    X_LUT4 C18832(
      .ADR0 (VCC),
      .ADR1 (\bridge/in_reg_cbe_out [1]),
      .ADR2 (syn16992),
      .ADR3 (VCC),
      .O (\bridge/configuration/C285/N99/GROM )
    );
    defparam C18861.INIT = 16'h4444;
    X_LUT4 C18861(
      .ADR0 (\bridge/in_reg_cbe_out [1]),
      .ADR1 (syn17097),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/configuration/C285/N99/FROM )
    );
    X_BUF \bridge/configuration/C285/N99/YUSED (
      .I (\bridge/configuration/C285/N99/GROM ),
      .O (\bridge/configuration/C280/N3 )
    );
    X_BUF \bridge/configuration/C285/N99/XUSED (
      .I (\bridge/configuration/C285/N99/FROM ),
      .O (\bridge/configuration/C285/N99 )
    );
    defparam C18824.INIT = 16'h0800;
    X_LUT4 C18824(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/configuration/C1925 ),
      .ADR2 (\bridge/in_reg_cbe_out [3]),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\bridge/configuration/C296/N24/GROM )
    );
    defparam C18843.INIT = 16'h0800;
    X_LUT4 C18843(
      .ADR0 (\bridge/configuration/C1953 ),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/in_reg_cbe_out [3]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C296/N24/FROM )
    );
    X_BUF \bridge/configuration/C296/N24/YUSED (
      .I (\bridge/configuration/C296/N24/GROM ),
      .O (\bridge/configuration/C301/N3 )
    );
    X_BUF \bridge/configuration/C296/N24/XUSED (
      .I (\bridge/configuration/C296/N24/FROM ),
      .O (\bridge/configuration/C296/N24 )
    );
    defparam C18808.INIT = 16'h4000;
    X_LUT4 C18808(
      .ADR0 (\bridge/in_reg_cbe_out [0]),
      .ADR1 (syn16934),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/configuration/C2240 ),
      .O (\bridge/configuration/C293/N14/GROM )
    );
    defparam C18812.INIT = 16'h4000;
    X_LUT4 C18812(
      .ADR0 (\bridge/in_reg_cbe_out [0]),
      .ADR1 (\bridge/configuration/C1959 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C293/N14/FROM )
    );
    X_BUF \bridge/configuration/C293/N14/YUSED (
      .I (\bridge/configuration/C293/N14/GROM ),
      .O (\bridge/configuration/C288/N39 )
    );
    X_BUF \bridge/configuration/C293/N14/XUSED (
      .I (\bridge/configuration/C293/N14/FROM ),
      .O (\bridge/configuration/C293/N14 )
    );
    defparam C18576.INIT = 16'hEAC0;
    X_LUT4 C18576(
      .ADR0 (syn136386),
      .ADR1 (syn136384),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [13]),
      .ADR3 (\bridge/pci_target_unit/fifos_pcir_data_out [13]),
      .O (\syn180261/GROM )
    );
    defparam C18621.INIT = 16'hECA0;
    X_LUT4 C18621(
      .ADR0 (syn136386),
      .ADR1 (syn136384),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [10]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [10]),
      .O (\syn180261/FROM )
    );
    X_BUF \syn180261/YUSED (
      .I (\syn180261/GROM ),
      .O (syn180385)
    );
    X_BUF \syn180261/XUSED (
      .I (\syn180261/FROM ),
      .O (syn180261)
    );
    defparam C18568.INIT = 16'hF888;
    X_LUT4 C18568(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [14]),
      .ADR2 (syn17068),
      .ADR3 (syn60110),
      .O (\bridge/configuration/C286/N19/GROM )
    );
    defparam C18906.INIT = 16'h0A00;
    X_LUT4 C18906(
      .ADR0 (syn60110),
      .ADR1 (VCC),
      .ADR2 (\bridge/in_reg_cbe_out [3]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C286/N19/FROM )
    );
    X_BUF \bridge/configuration/C286/N19/YUSED (
      .I (\bridge/configuration/C286/N19/GROM ),
      .O (syn180416)
    );
    X_BUF \bridge/configuration/C286/N19/XUSED (
      .I (\bridge/configuration/C286/N19/FROM ),
      .O (\bridge/configuration/C286/N19 )
    );
    defparam C17960.INIT = 16'h8421;
    X_LUT4 C17960(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [21]),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [20]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[21]/GROM )
    );
    defparam C19374.INIT = 16'hFFAA;
    X_LUT4 C19374(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[21]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<21>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[21]/GROM ),
      .O (syn181993)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<21>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[21]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [21])
    );
    defparam C17928.INIT = 16'h7BDE;
    X_LUT4 C17928(
      .ADR0 (\bridge/pci_target_unit/fifos/outGreyCount [2]),
      .ADR1 (\bridge/pci_target_unit/fifos/outGreyCount [3]),
      .ADR2 (\bridge/pci_target_unit/fifos/inGreyCount [2]),
      .ADR3 (\bridge/pci_target_unit/fifos/inGreyCount [3]),
      .O (\syn182037/GROM )
    );
    X_BUF \syn182037/YUSED (
      .I (\syn182037/GROM ),
      .O (syn182037)
    );
    defparam C17792.INIT = 16'hB000;
    X_LUT4 C17792(
      .ADR0 (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .ADR1 (\bridge/pci_target_unit/del_sync/req_comp_pending ),
      .ADR2 (syn19366),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/rd_request ),
      .O (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/GROM )
    );
    defparam C19308.INIT = 16'h00F0;
    X_LUT4 C19308(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/req_comp_pending ),
      .ADR3 (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .O (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/FROM )
    );
    X_INV \bridge/pci_target_unit/pci_target_sm/read_completed_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/read_completed_reg/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/GROM ),
      .O (syn182355)
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/read_completed_reg/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_read_completed_out )
    );
    X_FF \bridge/pci_target_unit/pci_target_sm/read_completed_reg_reg (
      .I (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_sm/read_completed_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_sm/read_completed_reg/FFX/ASYNC_FF_GSR_OR_146 (
      .I0 (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_sm/read_completed_reg/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C19705.INIT = 16'hECA0;
    X_LUT4 C19705(
      .ADR0 (\bridge/configuration/wb_addr_mask1 [18]),
      .ADR1 (\bridge/configuration/C2370 ),
      .ADR2 (\bridge/configuration/C2320 ),
      .ADR3 (\bridge/configuration/pci_base_addr0 [18]),
      .O (\syn177990/GROM )
    );
    defparam C19718.INIT = 16'hEAC0;
    X_LUT4 C19718(
      .ADR0 (\bridge/configuration/C2370 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [19]),
      .ADR2 (\bridge/configuration/C2320 ),
      .ADR3 (\bridge/configuration/pci_base_addr0 [19]),
      .O (\syn177990/FROM )
    );
    X_BUF \syn177990/YUSED (
      .I (\syn177990/GROM ),
      .O (syn178023)
    );
    X_BUF \syn177990/XUSED (
      .I (\syn177990/FROM ),
      .O (syn177990)
    );
    defparam C19553.INIT = 16'hFCCC;
    X_LUT4 C19553(
      .ADR0 (VCC),
      .ADR1 (syn24326),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [6]),
      .ADR3 (syn17745),
      .O (\syn24470/GROM )
    );
    defparam C19573.INIT = 16'hEAEA;
    X_LUT4 C19573(
      .ADR0 (syn24326),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [8]),
      .ADR2 (syn17745),
      .ADR3 (VCC),
      .O (\syn24470/FROM )
    );
    X_BUF \syn24470/YUSED (
      .I (\syn24470/GROM ),
      .O (syn24472)
    );
    X_BUF \syn24470/XUSED (
      .I (\syn24470/FROM ),
      .O (syn24470)
    );
    defparam C19377.INIT = 16'hFAFA;
    X_LUT4 C19377(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[24]/GROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<24>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[24]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [24])
    );
    defparam C18825.INIT = 16'h0800;
    X_LUT4 C18825(
      .ADR0 (\bridge/configuration/C1955 ),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/in_reg_cbe_out [0]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C298/N3/GROM )
    );
    defparam C18842.INIT = 16'h0080;
    X_LUT4 C18842(
      .ADR0 (\bridge/configuration/C1941 ),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/in_reg_cbe_out [0]),
      .O (\bridge/configuration/C298/N3/FROM )
    );
    X_BUF \bridge/configuration/C298/N3/YUSED (
      .I (\bridge/configuration/C298/N3/GROM ),
      .O (\bridge/configuration/C295/N3 )
    );
    X_BUF \bridge/configuration/C298/N3/XUSED (
      .I (\bridge/configuration/C298/N3/FROM ),
      .O (\bridge/configuration/C298/N3 )
    );
    defparam C18809.INIT = 16'h8000;
    X_LUT4 C18809(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (\bridge/pciu_conf_offset_out [5]),
      .ADR3 (\bridge/pciu_conf_offset_out [4]),
      .O (\syn179762/GROM )
    );
    defparam C18835.INIT = 16'hAABF;
    X_LUT4 C18835(
      .ADR0 (\bridge/pciu_conf_offset_out [5]),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (\bridge/pciu_conf_offset_out [2]),
      .ADR3 (\bridge/pciu_conf_offset_out [4]),
      .O (\syn179762/FROM )
    );
    X_BUF \syn179762/YUSED (
      .I (\syn179762/GROM ),
      .O (\bridge/configuration/C2240 )
    );
    X_BUF \syn179762/XUSED (
      .I (\syn179762/FROM ),
      .O (syn179762)
    );
    defparam C18745.INIT = 16'hF888;
    X_LUT4 C18745(
      .ADR0 (\bridge/configuration/C1929 ),
      .ADR1 (\bridge/configuration/config_addr[2] ),
      .ADR2 (\bridge/configuration/perr_int_en ),
      .ADR3 (\bridge/configuration/C1925 ),
      .O (\syn178462/GROM )
    );
    defparam C19514.INIT = 16'hF888;
    X_LUT4 C19514(
      .ADR0 (\bridge/configuration/C2304 ),
      .ADR1 (\bridge/configuration/wb_err_addr [2]),
      .ADR2 (\bridge/configuration/C2296 ),
      .ADR3 (\bridge/configuration/config_addr[2] ),
      .O (\syn178462/FROM )
    );
    X_BUF \syn178462/YUSED (
      .I (\syn178462/GROM ),
      .O (syn179949)
    );
    X_BUF \syn178462/XUSED (
      .I (\syn178462/FROM ),
      .O (syn178462)
    );
    defparam C18737.INIT = 16'hC088;
    X_LUT4 C18737(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [2]),
      .ADR1 (syn19366),
      .ADR2 (\bridge/pci_target_unit/fifos_pcir_data_out [2]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_291/cell0 ),
      .O (\syn178883/GROM )
    );
    defparam C19311.INIT = 16'h4000;
    X_LUT4 C19311(
      .ADR0 (\bridge/pci_target_unit/fifos_pciw_full_out ),
      .ADR1 (syn19366),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/wr_to_fifo ),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .O (\syn178883/FROM )
    );
    X_BUF \syn178883/YUSED (
      .I (\syn178883/GROM ),
      .O (syn179957)
    );
    X_BUF \syn178883/XUSED (
      .I (\syn178883/FROM ),
      .O (syn178883)
    );
    defparam C18585.INIT = 16'hF888;
    X_LUT4 C18585(
      .ADR0 (\bridge/configuration/config_addr[13] ),
      .ADR1 (\bridge/configuration/C1929 ),
      .ADR2 (\bridge/configuration/wb_err_data [13]),
      .ADR3 (\bridge/configuration/C1935 ),
      .O (\syn180316/GROM )
    );
    defparam C18603.INIT = 16'hEAC0;
    X_LUT4 C18603(
      .ADR0 (\bridge/configuration/config_addr[12] ),
      .ADR1 (\bridge/configuration/C1935 ),
      .ADR2 (\bridge/configuration/wb_err_data [12]),
      .ADR3 (\bridge/configuration/C1929 ),
      .O (\syn180316/FROM )
    );
    X_BUF \syn180316/YUSED (
      .I (\syn180316/GROM ),
      .O (syn180368)
    );
    X_BUF \syn180316/XUSED (
      .I (\syn180316/FROM ),
      .O (syn180316)
    );
    defparam C18569.INIT = 16'hECCC;
    X_LUT4 C18569(
      .ADR0 (syn17005),
      .ADR1 (\bridge/configuration/C2001 ),
      .ADR2 (syn17004),
      .ADR3 (syn179659),
      .O (\syn17120/GROM )
    );
    defparam C18779.INIT = 16'h8000;
    X_LUT4 C18779(
      .ADR0 (syn16914),
      .ADR1 (syn60111),
      .ADR2 (syn17005),
      .ADR3 (syn179659),
      .O (\syn17120/FROM )
    );
    X_BUF \syn17120/YUSED (
      .I (\syn17120/GROM ),
      .O (syn48754)
    );
    X_BUF \syn17120/XUSED (
      .I (\syn17120/FROM ),
      .O (syn17120)
    );
    defparam C18497.INIT = 16'hF888;
    X_LUT4 C18497(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [18]),
      .ADR1 (syn20493),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [18]),
      .O (\syn180270/GROM )
    );
    defparam C18612.INIT = 16'hEAC0;
    X_LUT4 C18612(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [11]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [11]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .ADR3 (syn20493),
      .O (\syn180270/FROM )
    );
    X_BUF \syn180270/YUSED (
      .I (\syn180270/GROM ),
      .O (syn180623)
    );
    X_BUF \syn180270/XUSED (
      .I (\syn180270/FROM ),
      .O (syn180270)
    );
    defparam C17961.INIT = 16'h9009;
    X_LUT4 C17961(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [23]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [22]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[23]/GROM )
    );
    defparam C19376.INIT = 16'hFAFA;
    X_LUT4 C19376(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[23]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<23>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[23]/GROM ),
      .O (syn181992)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<23>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[23]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [23])
    );
    defparam C17785.INIT = 16'hFAFF;
    X_LUT4 C17785(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/S_198/cell0 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_cycle_count [16]),
      .ADR3 (\bridge/pci_target_unit/del_sync/req_comp_pending_sample ),
      .O (\N12541/GROM )
    );
    defparam C17788.INIT = 16'hFFBB;
    X_LUT4 C17788(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/S_198/cell0 ),
      .ADR1 (\bridge/pci_target_unit/del_sync/req_done_reg ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/comp_cycle_count [16]),
      .O (\N12541/FROM )
    );
    X_BUF \N12541/YUSED (
      .I (\N12541/GROM ),
      .O (N12540)
    );
    X_BUF \N12541/XUSED (
      .I (\N12541/FROM ),
      .O (N12541)
    );
    defparam \bridge/pci_target_unit/del_sync/req_rty_exp_reg/F .INIT = 16'h0000;
    X_LUT4 \bridge/pci_target_unit/del_sync/req_rty_exp_reg/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_reg/FROM )
    );
    X_INV \bridge/pci_target_unit/del_sync/req_rty_exp_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_reg/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/del_sync/req_rty_exp_reg/XUSED (
      .I (\bridge/pci_target_unit/del_sync/req_rty_exp_reg/FROM ),
      .O (GLOBAL_LOGIC0_0)
    );
    X_FF \bridge/pci_target_unit/del_sync/req_rty_exp_reg_reg (
      .I (\bridge/pci_target_unit/del_sync/sync_req_rty_exp ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/req_rty_exp_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_reg )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/req_rty_exp_reg/FFY/ASYNC_FF_GSR_OR_147 (
      .I0 (\bridge/pci_target_unit/del_sync/req_rty_exp_reg/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync/req_rty_exp_reg/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/sync_req_rty_exp ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg/FFY/ASYNC_FF_GSR_OR_148 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/req_rty_exp_reg/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19706.INIT = 16'hEAC0;
    X_LUT4 C19706(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [18]),
      .ADR1 (\bridge/configuration/pci_err_addr [18]),
      .ADR2 (\bridge/configuration/C2338 ),
      .ADR3 (\bridge/configuration/C2318 ),
      .O (\syn177989/GROM )
    );
    defparam C19719.INIT = 16'hECA0;
    X_LUT4 C19719(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [19]),
      .ADR2 (\bridge/configuration/pci_err_addr [19]),
      .ADR3 (\bridge/configuration/C2318 ),
      .O (\syn177989/FROM )
    );
    X_BUF \syn177989/YUSED (
      .I (\syn177989/GROM ),
      .O (syn178022)
    );
    X_BUF \syn177989/XUSED (
      .I (\syn177989/FROM ),
      .O (syn177989)
    );
    defparam C19490.INIT = 16'hEAC0;
    X_LUT4 C19490(
      .ADR0 (\bridge/conf_pci_mem_io1_out ),
      .ADR1 (\bridge/conf_io_space_enable_out ),
      .ADR2 (syn24559),
      .ADR3 (syn16928),
      .O (\syn177710/GROM )
    );
    defparam C19835.INIT = 16'hF888;
    X_LUT4 C19835(
      .ADR0 (\bridge/configuration/status_bit15_11 [11]),
      .ADR1 (syn24559),
      .ADR2 (syn16928),
      .ADR3 (syn17054),
      .O (\syn177710/FROM )
    );
    X_BUF \syn177710/YUSED (
      .I (\syn177710/GROM ),
      .O (syn178528)
    );
    X_BUF \syn177710/XUSED (
      .I (\syn177710/FROM ),
      .O (syn177710)
    );
    defparam C18850.INIT = 16'h0080;
    X_LUT4 C18850(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/configuration/C1989 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/in_reg_cbe_out [3]),
      .O (\bridge/configuration/C294/N29/GROM )
    );
    defparam C18899.INIT = 16'h0080;
    X_LUT4 C18899(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1955 ),
      .ADR3 (\bridge/in_reg_cbe_out [3]),
      .O (\bridge/configuration/C294/N29/FROM )
    );
    X_BUF \bridge/configuration/C294/N29/YUSED (
      .I (\bridge/configuration/C294/N29/GROM ),
      .O (\bridge/configuration/C290/N3 )
    );
    X_BUF \bridge/configuration/C294/N29/XUSED (
      .I (\bridge/configuration/C294/N29/FROM ),
      .O (\bridge/configuration/C294/N29 )
    );
    defparam C18586.INIT = 16'hECA0;
    X_LUT4 C18586(
      .ADR0 (\bridge/configuration/pci_base_addr0 [13]),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [13]),
      .ADR2 (\bridge/configuration/C2003 ),
      .ADR3 (\bridge/configuration/C1989 ),
      .O (\syn180315/GROM )
    );
    defparam C18604.INIT = 16'hF888;
    X_LUT4 C18604(
      .ADR0 (\bridge/configuration/C1989 ),
      .ADR1 (\bridge/configuration/pci_addr_mask1 [12]),
      .ADR2 (\bridge/configuration/C2003 ),
      .ADR3 (\bridge/configuration/pci_base_addr0 [12]),
      .O (\syn180315/FROM )
    );
    X_BUF \syn180315/YUSED (
      .I (\syn180315/GROM ),
      .O (syn180367)
    );
    X_BUF \syn180315/XUSED (
      .I (\syn180315/FROM ),
      .O (syn180315)
    );
    defparam C17954.INIT = 16'h8421;
    X_LUT4 C17954(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [10]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [11]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [10]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [11]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[11]/GROM )
    );
    defparam C19340.INIT = 16'hFFF0;
    X_LUT4 C19340(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [11]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[11]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<11>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[11]/GROM ),
      .O (syn181998)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<11>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[11]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [11])
    );
    defparam C19731.INIT = 16'hF888;
    X_LUT4 C19731(
      .ADR0 (\bridge/configuration/C2302 ),
      .ADR1 (\bridge/configuration/wb_err_data [20]),
      .ADR2 (\bridge/configuration/C2318 ),
      .ADR3 (\bridge/configuration/wb_tran_addr1 [20]),
      .O (\syn177922/GROM )
    );
    defparam C19744.INIT = 16'hECA0;
    X_LUT4 C19744(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [21]),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (\bridge/configuration/C2318 ),
      .ADR3 (\bridge/configuration/wb_err_data [21]),
      .O (\syn177922/FROM )
    );
    X_BUF \syn177922/YUSED (
      .I (\syn177922/GROM ),
      .O (syn177955)
    );
    X_BUF \syn177922/XUSED (
      .I (\syn177922/FROM ),
      .O (syn177922)
    );
    defparam C19619.INIT = 16'hECA0;
    X_LUT4 C19619(
      .ADR0 (\bridge/configuration/pci_base_addr0 [12]),
      .ADR1 (\bridge/configuration/pci_err_addr [12]),
      .ADR2 (\bridge/configuration/C2370 ),
      .ADR3 (\bridge/configuration/C2338 ),
      .O (\syn178094/GROM )
    );
    defparam C19678.INIT = 16'hECA0;
    X_LUT4 C19678(
      .ADR0 (\bridge/configuration/pci_err_addr [16]),
      .ADR1 (\bridge/configuration/pci_base_addr0 [16]),
      .ADR2 (\bridge/configuration/C2338 ),
      .ADR3 (\bridge/configuration/C2370 ),
      .O (\syn178094/FROM )
    );
    X_BUF \syn178094/YUSED (
      .I (\syn178094/GROM ),
      .O (syn178238)
    );
    X_BUF \syn178094/XUSED (
      .I (\syn178094/FROM ),
      .O (syn178094)
    );
    defparam C19547.INIT = 16'hEAC0;
    X_LUT4 C19547(
      .ADR0 (\bridge/configuration/config_addr[6] ),
      .ADR1 (\bridge/configuration/pci_err_addr [6]),
      .ADR2 (syn16984),
      .ADR3 (syn17079),
      .O (\syn178311/GROM )
    );
    defparam C19576.INIT = 16'hEAC0;
    X_LUT4 C19576(
      .ADR0 (\bridge/configuration/config_addr[9] ),
      .ADR1 (syn17078),
      .ADR2 (\bridge/configuration/wb_err_addr [9]),
      .ADR3 (syn17079),
      .O (\syn178311/FROM )
    );
    X_BUF \syn178311/YUSED (
      .I (\syn178311/GROM ),
      .O (syn178373)
    );
    X_BUF \syn178311/XUSED (
      .I (\syn178311/FROM ),
      .O (syn178311)
    );
    defparam C18819.INIT = 16'h80C0;
    X_LUT4 C18819(
      .ADR0 (ERR_I),
      .ADR1 (\bridge/configuration/pci_error_en ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR3 (ACK_I),
      .O (\syn179789/GROM )
    );
    X_BUF \syn179789/YUSED (
      .I (\syn179789/GROM ),
      .O (syn179789)
    );
    defparam C18587.INIT = 16'hECA0;
    X_LUT4 C18587(
      .ADR0 (\bridge/configuration/C1987 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [13]),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [13]),
      .ADR3 (\bridge/configuration/C1951 ),
      .O (\syn180314/GROM )
    );
    defparam C18605.INIT = 16'hEAC0;
    X_LUT4 C18605(
      .ADR0 (\bridge/configuration/C1987 ),
      .ADR1 (\bridge/configuration/C1951 ),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [12]),
      .ADR3 (\bridge/configuration/pci_tran_addr1 [12]),
      .O (\syn180314/FROM )
    );
    X_BUF \syn180314/YUSED (
      .I (\syn180314/GROM ),
      .O (syn180366)
    );
    X_BUF \syn180314/XUSED (
      .I (\syn180314/FROM ),
      .O (syn180314)
    );
    defparam C17947.INIT = 16'h8421;
    X_LUT4 C17947(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [26]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [27]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[27]/GROM )
    );
    defparam C19380.INIT = 16'hFFF0;
    X_LUT4 C19380(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[27]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<27>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[27]/GROM ),
      .O (syn181990)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<27>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[27]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [27])
    );
    defparam C19572.INIT = 16'h8080;
    X_LUT4 C19572(
      .ADR0 (\bridge/configuration/C2302 ),
      .ADR1 (\bridge/configuration/wb_err_data [8]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR3 (VCC),
      .O (\syn17077/GROM )
    );
    defparam C19592.INIT = 16'hC0C0;
    X_LUT4 C19592(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR2 (\bridge/configuration/C2334 ),
      .ADR3 (VCC),
      .O (\syn17077/FROM )
    );
    X_BUF \syn17077/YUSED (
      .I (\syn17077/GROM ),
      .O (syn18636)
    );
    X_BUF \syn17077/XUSED (
      .I (\syn17077/FROM ),
      .O (syn17077)
    );
    defparam C18908.INIT = 16'h0044;
    X_LUT4 C18908(
      .ADR0 (\bridge/in_reg_cbe_out [3]),
      .ADR1 (\bridge/configuration/C2003 ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[3]/GROM )
    );
    defparam C19215.INIT = 16'hDD88;
    X_LUT4 C19215(
      .ADR0 (\bridge/pci_target_unit/pcit_sm_rdy_out ),
      .ADR1 (\bridge/pci_target_unit/pcit_if_bc_out [3]),
      .ADR2 (VCC),
      .ADR3 (\bridge/in_reg_cbe_out [3]),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[3]/FROM )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out<3>/YUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[3]/GROM ),
      .O (\bridge/configuration/C338/N3 )
    );
    X_BUF \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out<3>/XUSED (
      .I (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out[3]/FROM ),
      .O (\bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out [3])
    );
    defparam C18852.INIT = 16'h0080;
    X_LUT4 C18852(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR2 (\bridge/configuration/C1987 ),
      .ADR3 (\bridge/in_reg_cbe_out [1]),
      .O (\bridge/configuration/C290/N99/GROM )
    );
    defparam C18855.INIT = 16'h0080;
    X_LUT4 C18855(
      .ADR0 (\bridge/configuration/C1989 ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/in_reg_cbe_out [1]),
      .O (\bridge/configuration/C290/N99/FROM )
    );
    X_BUF \bridge/configuration/C290/N99/YUSED (
      .I (\bridge/configuration/C290/N99/GROM ),
      .O (\bridge/configuration/C291/N94 )
    );
    X_BUF \bridge/configuration/C290/N99/XUSED (
      .I (\bridge/configuration/C290/N99/FROM ),
      .O (\bridge/configuration/C290/N99 )
    );
    defparam C18596.INIT = 16'hC888;
    X_LUT4 C18596(
      .ADR0 (syn120382),
      .ADR1 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR2 (syn17070),
      .ADR3 (syn16927),
      .O (\syn21466/GROM )
    );
    defparam C18348.INIT = 16'h8000;
    X_LUT4 C18348(
      .ADR0 (\bridge/out_bckp_tar_ad_en_out ),
      .ADR1 (\bridge/conf_pci_am1_out [15]),
      .ADR2 (syn16927),
      .ADR3 (\bridge/conf_pci_ba1_out [15]),
      .O (\syn21466/FROM )
    );
    X_BUF \syn21466/YUSED (
      .I (\syn21466/GROM ),
      .O (syn180336)
    );
    X_BUF \syn21466/XUSED (
      .I (\syn21466/FROM ),
      .O (syn21466)
    );
    defparam C17956.INIT = 16'h8241;
    X_LUT4 C17956(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [15]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [14]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[15]/GROM )
    );
    defparam C19344.INIT = 16'hEEEE;
    X_LUT4 C19344(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[15]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<15>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[15]/GROM ),
      .O (syn181996)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<15>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[15]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [15])
    );
    defparam C17948.INIT = 16'h8241;
    X_LUT4 C17948(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [29]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [28]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[29]/GROM )
    );
    defparam C19382.INIT = 16'hFCFC;
    X_LUT4 C19382(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[29]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<29>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[29]/GROM ),
      .O (syn181989)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<29>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[29]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [29])
    );
    defparam C19805.INIT = 16'hAA00;
    X_LUT4 C19805(
      .ADR0 (\bridge/conf_pci_am1_out [13]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_pci_ba1_out [13]),
      .O (\syn17056/GROM )
    );
    X_BUF \syn17056/YUSED (
      .I (\syn17056/GROM ),
      .O (syn17056)
    );
    defparam C19725.INIT = 16'hECA0;
    X_LUT4 C19725(
      .ADR0 (\bridge/configuration/C2296 ),
      .ADR1 (\bridge/configuration/wb_err_addr [20]),
      .ADR2 (\bridge/configuration/config_addr[20] ),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn177925/GROM )
    );
    defparam C19738.INIT = 16'hF888;
    X_LUT4 C19738(
      .ADR0 (\bridge/configuration/config_addr[21] ),
      .ADR1 (\bridge/configuration/C2296 ),
      .ADR2 (\bridge/configuration/wb_err_addr [21]),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn177925/FROM )
    );
    X_BUF \syn177925/YUSED (
      .I (\syn177925/GROM ),
      .O (syn177958)
    );
    X_BUF \syn177925/XUSED (
      .I (\syn177925/FROM ),
      .O (syn177925)
    );
    defparam C19709.INIT = 16'hF888;
    X_LUT4 C19709(
      .ADR0 (\bridge/configuration/pci_base_addr0 [19]),
      .ADR1 (syn16930),
      .ADR2 (syn17745),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [19]),
      .O (\syn177869/GROM )
    );
    defparam C19761.INIT = 16'hECA0;
    X_LUT4 C19761(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [23]),
      .ADR1 (\bridge/configuration/pci_base_addr0 [23]),
      .ADR2 (syn17745),
      .ADR3 (syn16930),
      .O (\syn177869/FROM )
    );
    X_BUF \syn177869/YUSED (
      .I (\syn177869/GROM ),
      .O (syn178002)
    );
    X_BUF \syn177869/XUSED (
      .I (\syn177869/FROM ),
      .O (syn177869)
    );
    defparam C19629.INIT = 16'hC000;
    X_LUT4 C19629(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_base_addr1 [13]),
      .ADR2 (\bridge/configuration/pci_addr_mask1 [13]),
      .ADR3 (\bridge/configuration/C2360 ),
      .O (\syn18087/GROM )
    );
    defparam C19788.INIT = 16'h8080;
    X_LUT4 C19788(
      .ADR0 (\bridge/configuration/C2360 ),
      .ADR1 (\bridge/conf_pci_ba1_out [12]),
      .ADR2 (\bridge/conf_pci_am1_out [12]),
      .ADR3 (VCC),
      .O (\syn18087/FROM )
    );
    X_BUF \syn18087/YUSED (
      .I (\syn18087/GROM ),
      .O (syn18491)
    );
    X_BUF \syn18087/XUSED (
      .I (\syn18087/FROM ),
      .O (syn18087)
    );
    defparam C19581.INIT = 16'hFAAA;
    X_LUT4 C19581(
      .ADR0 (syn24326),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [9]),
      .ADR3 (syn17745),
      .O (\syn24466/GROM )
    );
    defparam C19597.INIT = 16'hEAEA;
    X_LUT4 C19597(
      .ADR0 (syn24326),
      .ADR1 (syn17745),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [10]),
      .ADR3 (VCC),
      .O (\syn24466/FROM )
    );
    X_BUF \syn24466/YUSED (
      .I (\syn24466/GROM ),
      .O (syn24468)
    );
    X_BUF \syn24466/XUSED (
      .I (\syn24466/FROM ),
      .O (syn24466)
    );
    defparam C19493.INIT = 16'hF888;
    X_LUT4 C19493(
      .ADR0 (\bridge/configuration/C2322 ),
      .ADR1 (\bridge/conf_wb_mem_io1_out ),
      .ADR2 (\bridge/configuration/pci_err_addr [0]),
      .ADR3 (\bridge/configuration/C2338 ),
      .O (\syn16984/GROM )
    );
    defparam C19588.INIT = 16'hAA00;
    X_LUT4 C19588(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C2338 ),
      .O (\syn16984/FROM )
    );
    X_BUF \syn16984/YUSED (
      .I (\syn16984/GROM ),
      .O (syn178516)
    );
    X_BUF \syn16984/XUSED (
      .I (\syn16984/FROM ),
      .O (syn16984)
    );
    defparam C19485.INIT = 16'h0033;
    X_LUT4 C19485(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .O (\syn178535/GROM )
    );
    defparam \syn178535/F .INIT = 16'h0000;
    X_LUT4 \syn178535/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn178535/FROM )
    );
    X_BUF \syn178535/YUSED (
      .I (\syn178535/GROM ),
      .O (syn178535)
    );
    X_BUF \syn178535/XUSED (
      .I (\syn178535/FROM ),
      .O (GLOBAL_LOGIC0)
    );
    defparam C18853.INIT = 16'h0080;
    X_LUT4 C18853(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1987 ),
      .ADR3 (\bridge/in_reg_cbe_out [2]),
      .O (\bridge/configuration/C296/N64/GROM )
    );
    defparam C18854.INIT = 16'h0080;
    X_LUT4 C18854(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/in_reg_cbe_out [2]),
      .O (\bridge/configuration/C296/N64/FROM )
    );
    X_BUF \bridge/configuration/C296/N64/YUSED (
      .I (\bridge/configuration/C296/N64/GROM ),
      .O (\bridge/configuration/C291/N59 )
    );
    X_BUF \bridge/configuration/C296/N64/XUSED (
      .I (\bridge/configuration/C296/N64/FROM ),
      .O (\bridge/configuration/C296/N64 )
    );
    defparam C18845.INIT = 16'h0080;
    X_LUT4 C18845(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR2 (\bridge/configuration/C1953 ),
      .ADR3 (\bridge/in_reg_cbe_out [1]),
      .O (\bridge/configuration/C297/N84/GROM )
    );
    defparam C18847.INIT = 16'h4000;
    X_LUT4 C18847(
      .ADR0 (\bridge/in_reg_cbe_out [1]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/configuration/C1951 ),
      .O (\bridge/configuration/C297/N84/FROM )
    );
    X_BUF \bridge/configuration/C297/N84/YUSED (
      .I (\bridge/configuration/C297/N84/GROM ),
      .O (\bridge/configuration/C296/N89 )
    );
    X_BUF \bridge/configuration/C297/N84/XUSED (
      .I (\bridge/configuration/C297/N84/FROM ),
      .O (\bridge/configuration/C297/N84 )
    );
    defparam C18829.INIT = 16'h4180;
    X_LUT4 C18829(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [4]),
      .ADR2 (\bridge/pciu_conf_offset_out [7]),
      .ADR3 (\bridge/pciu_conf_offset_out [5]),
      .O (\syn179761/GROM )
    );
    defparam C18836.INIT = 16'h3322;
    X_LUT4 C18836(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [5]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pciu_conf_offset_out [4]),
      .O (\syn179761/FROM )
    );
    X_BUF \syn179761/YUSED (
      .I (\syn179761/GROM ),
      .O (syn179776)
    );
    X_BUF \syn179761/XUSED (
      .I (\syn179761/FROM ),
      .O (syn179761)
    );
    defparam C18757.INIT = 16'hF888;
    X_LUT4 C18757(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (\bridge/configuration/wb_err_data [1]),
      .ADR2 (\bridge/configuration/C1925 ),
      .ADR3 (\bridge/configuration/error_int_en ),
      .O (\syn179847/GROM )
    );
    defparam C18793.INIT = 16'hEAC0;
    X_LUT4 C18793(
      .ADR0 (\bridge/configuration/C1935 ),
      .ADR1 (\bridge/configuration/config_addr[0] ),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/configuration/wb_err_data [0]),
      .O (\syn179847/FROM )
    );
    X_BUF \syn179847/YUSED (
      .I (\syn179847/GROM ),
      .O (syn179911)
    );
    X_BUF \syn179847/XUSED (
      .I (\syn179847/FROM ),
      .O (syn179847)
    );
    defparam C18749.INIT = 16'hECA0;
    X_LUT4 C18749(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_data_out [1]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_next_data_out [1]),
      .ADR2 (syn20493),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/N147 ),
      .O (\syn179894/GROM )
    );
    X_BUF \syn179894/YUSED (
      .I (\syn179894/GROM ),
      .O (syn179894)
    );
    defparam C18685.INIT = 16'hEAC0;
    X_LUT4 C18685(
      .ADR0 (syn17014),
      .ADR1 (syn17015),
      .ADR2 (\bridge/configuration/wb_err_data [6]),
      .ADR3 (\bridge/configuration/wb_err_addr [6]),
      .O (\syn180052/GROM )
    );
    defparam C18699.INIT = 16'hEAC0;
    X_LUT4 C18699(
      .ADR0 (syn17014),
      .ADR1 (syn17015),
      .ADR2 (\bridge/configuration/wb_err_data [5]),
      .ADR3 (\bridge/configuration/wb_err_addr [5]),
      .O (\syn180052/FROM )
    );
    X_BUF \syn180052/YUSED (
      .I (\syn180052/GROM ),
      .O (syn180083)
    );
    X_BUF \syn180052/XUSED (
      .I (\syn180052/FROM ),
      .O (syn180052)
    );
    defparam C17949.INIT = 16'h8421;
    X_LUT4 C17949(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .ADR1 (\bridge/pci_target_unit/del_sync_addr_out [30]),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [31]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[30]/GROM )
    );
    defparam C19383.INIT = 16'hFFAA;
    X_LUT4 C19383(
      .ADR0 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[30]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<30>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[30]/GROM ),
      .O (syn181988)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<30>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[30]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [30])
    );
    defparam C17893.INIT = 16'h0400;
    X_LUT4 C17893(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_full_out ),
      .ADR1 (\bridge/pci_target_unit/del_sync_comp_req_pending_out ),
      .ADR2 (syn19577),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C81/N3 ),
      .O (\syn17020/GROM )
    );
    defparam C17903.INIT = 16'h0100;
    X_LUT4 C17903(
      .ADR0 (\bridge/pci_target_unit/fifos_pcir_full_out ),
      .ADR1 (\bridge/conf_pci_err_pending_out ),
      .ADR2 (syn19577),
      .ADR3 (\bridge/pci_target_unit/del_sync_comp_req_pending_out ),
      .O (\syn17020/FROM )
    );
    X_BUF \syn17020/YUSED (
      .I (\syn17020/GROM ),
      .O (syn16925)
    );
    X_BUF \syn17020/XUSED (
      .I (\syn17020/FROM ),
      .O (syn17020)
    );
    defparam C19654.INIT = 16'h8800;
    X_LUT4 C19654(
      .ADR0 (\bridge/configuration/pci_base_addr1 [15]),
      .ADR1 (syn16928),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/pci_addr_mask1 [15]),
      .O (\syn178035/GROM )
    );
    defparam C19696.INIT = 16'hEAC0;
    X_LUT4 C19696(
      .ADR0 (syn17063),
      .ADR1 (syn17745),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [18]),
      .ADR3 (syn16928),
      .O (\syn178035/FROM )
    );
    X_BUF \syn178035/YUSED (
      .I (\syn178035/GROM ),
      .O (syn18431)
    );
    X_BUF \syn178035/XUSED (
      .I (\syn178035/FROM ),
      .O (syn178035)
    );
    defparam C19494.INIT = 16'hF000;
    X_LUT4 C19494(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/C2296 ),
      .ADR3 (\bridge/configuration/config_addr[0] ),
      .O (\syn178240/GROM )
    );
    defparam C19614.INIT = 16'hEAC0;
    X_LUT4 C19614(
      .ADR0 (\bridge/configuration/C2304 ),
      .ADR1 (\bridge/configuration/config_addr[12] ),
      .ADR2 (\bridge/configuration/C2296 ),
      .ADR3 (\bridge/configuration/wb_err_addr [12]),
      .O (\syn178240/FROM )
    );
    X_BUF \syn178240/YUSED (
      .I (\syn178240/GROM ),
      .O (syn178517)
    );
    X_BUF \syn178240/XUSED (
      .I (\syn178240/FROM ),
      .O (syn178240)
    );
    defparam C19398.INIT = 16'h0005;
    X_LUT4 C19398(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_last ),
      .ADR1 (VCC),
      .ADR2 (\bridge/in_reg_trdy_out ),
      .ADR3 (\bridge/in_reg_devsel_out ),
      .O (\syn19064/GROM )
    );
    defparam C19410.INIT = 16'hDDD0;
    X_LUT4 C19410(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort1 ),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/mabort2 ),
      .ADR2 (\bridge/in_reg_trdy_out ),
      .ADR3 (\bridge/in_reg_devsel_out ),
      .O (\syn19064/FROM )
    );
    X_BUF \syn19064/YUSED (
      .I (\syn19064/GROM ),
      .O (syn178711)
    );
    X_BUF \syn19064/XUSED (
      .I (\syn19064/FROM ),
      .O (syn19064)
    );
    defparam C18846.INIT = 16'h4000;
    X_LUT4 C18846(
      .ADR0 (\bridge/in_reg_cbe_out [3]),
      .ADR1 (\bridge/configuration/C1951 ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/pciu_conf_offset_out [8]),
      .O (\bridge/configuration/C291/N14/GROM )
    );
    defparam C18849.INIT = 16'h0080;
    X_LUT4 C18849(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR1 (\bridge/configuration/C1987 ),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/in_reg_cbe_out [3]),
      .O (\bridge/configuration/C291/N14/FROM )
    );
    X_BUF \bridge/configuration/C291/N14/YUSED (
      .I (\bridge/configuration/C291/N14/GROM ),
      .O (\bridge/configuration/C297/N29 )
    );
    X_BUF \bridge/configuration/C291/N14/XUSED (
      .I (\bridge/configuration/C291/N14/FROM ),
      .O (\bridge/configuration/C291/N14 )
    );
    defparam C18758.INIT = 16'hA000;
    X_LUT4 C18758(
      .ADR0 (\bridge/conf_pci_img_ctrl1_out [0]),
      .ADR1 (VCC),
      .ADR2 (syn60111),
      .ADR3 (syn60090),
      .O (\syn18784/GROM )
    );
    defparam C19508.INIT = 16'h8800;
    X_LUT4 C19508(
      .ADR0 (syn177632),
      .ADR1 (\bridge/conf_pci_img_ctrl1_out [0]),
      .ADR2 (VCC),
      .ADR3 (\bridge/configuration/C3488 ),
      .O (\syn18784/FROM )
    );
    X_BUF \syn18784/YUSED (
      .I (\syn18784/GROM ),
      .O (syn179910)
    );
    X_BUF \syn18784/XUSED (
      .I (\syn18784/FROM ),
      .O (syn18784)
    );
    defparam C18766.INIT = 16'hA000;
    X_LUT4 C18766(
      .ADR0 (syn16914),
      .ADR1 (VCC),
      .ADR2 (syn60111),
      .ADR3 (\bridge/configuration/C2268 ),
      .O (\syn179948/GROM )
    );
    defparam C18743.INIT = 16'hC000;
    X_LUT4 C18743(
      .ADR0 (VCC),
      .ADR1 (\bridge/configuration/pci_img_ctrl1 [2]),
      .ADR2 (syn60111),
      .ADR3 (syn60090),
      .O (\syn179948/FROM )
    );
    X_BUF \syn179948/YUSED (
      .I (\syn179948/GROM ),
      .O (syn17101)
    );
    X_BUF \syn179948/XUSED (
      .I (\syn179948/FROM ),
      .O (syn179948)
    );
    defparam C17798.INIT = 16'h2000;
    X_LUT4 C17798(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [2]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [3]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [1]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [0]),
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/GROM )
    );
    defparam C17800.INIT = 16'h6A00;
    X_LUT4 C17800(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [2]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [0]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [1]),
      .ADR3 (syn17006),
      .O (\bridge/pci_target_unit/wishbone_master/C103/N15 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<2>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/SRNOT )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<2>/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/GROM ),
      .O (syn23094)
    );
    X_FF \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt_reg<2> (
      .I (\bridge/pci_target_unit/wishbone_master/C103/N15 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/wishbone_master/C104/N6 ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt [2])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/wb_no_response_cnt<2>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/wb_no_response_cnt[2]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C19815.INIT = 16'hF888;
    X_LUT4 C19815(
      .ADR0 (\bridge/configuration/pci_err_data [26]),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (\bridge/configuration/pci_err_cs_bit31_24 [26]),
      .ADR3 (\bridge/configuration/C2340 ),
      .O (\syn177613/GROM )
    );
    defparam C19863.INIT = 16'hEAC0;
    X_LUT4 C19863(
      .ADR0 (\bridge/configuration/pci_err_cs_bit31_24 [29]),
      .ADR1 (\bridge/configuration/C2334 ),
      .ADR2 (\bridge/configuration/pci_err_data [29]),
      .ADR3 (\bridge/configuration/C2340 ),
      .O (\syn177613/FROM )
    );
    X_BUF \syn177613/YUSED (
      .I (\syn177613/GROM ),
      .O (syn177737)
    );
    X_BUF \syn177613/XUSED (
      .I (\syn177613/FROM ),
      .O (syn177613)
    );
    defparam C18863.INIT = 16'h2020;
    X_LUT4 C18863(
      .ADR0 (\bridge/out_bckp_devsel_out ),
      .ADR1 (\bridge/out_bckp_stop_out ),
      .ADR2 (\bridge/out_bckp_trdy_out ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy/GROM )
    );
    defparam C19138.INIT = 16'hCECC;
    X_LUT4 C19138(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/c_state [1]),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/stop_w_frm_irdy ),
      .ADR2 (\bridge/out_bckp_trdy_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/c_state [0]),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy/FROM )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy/YUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy/GROM ),
      .O (\bridge/pciu_pciif_tabort_set_out )
    );
    X_BUF \bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy/XUSED (
      .I (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy/FROM ),
      .O (\bridge/pci_target_unit/pci_target_sm/trdy_w_frm_irdy )
    );
    defparam C18687.INIT = 16'hECA0;
    X_LUT4 C18687(
      .ADR0 (syn17105),
      .ADR1 (\bridge/conf_cache_line_size_out [6]),
      .ADR2 (\bridge/configuration/interrupt_line [6]),
      .ADR3 (syn17102),
      .O (\syn178376/GROM )
    );
    defparam C19549.INIT = 16'hEAC0;
    X_LUT4 C19549(
      .ADR0 (\bridge/configuration/pci_err_data [6]),
      .ADR1 (\bridge/conf_cache_line_size_out [6]),
      .ADR2 (syn17081),
      .ADR3 (syn17077),
      .O (\syn178376/FROM )
    );
    X_BUF \syn178376/YUSED (
      .I (\syn178376/GROM ),
      .O (syn180081)
    );
    X_BUF \syn178376/XUSED (
      .I (\syn178376/FROM ),
      .O (syn178376)
    );
    defparam C17959.INIT = 16'h8421;
    X_LUT4 C17959(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .ADR2 (\bridge/pci_target_unit/del_sync_addr_out [18]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [19]),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[19]/GROM )
    );
    defparam C19372.INIT = 16'hEEEE;
    X_LUT4 C19372(
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out[19]/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<19>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[19]/GROM ),
      .O (syn181994)
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_sm_data_out<19>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_sm_data_out[19]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_sm_data_out [19])
    );
    defparam C19648.INIT = 16'hECA0;
    X_LUT4 C19648(
      .ADR0 (\bridge/configuration/C2370 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [14]),
      .ADR2 (\bridge/configuration/pci_base_addr0 [14]),
      .ADR3 (\bridge/configuration/C2320 ),
      .O (\syn178132/GROM )
    );
    defparam C19663.INIT = 16'hF888;
    X_LUT4 C19663(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [15]),
      .ADR2 (\bridge/configuration/C2370 ),
      .ADR3 (\bridge/configuration/pci_base_addr0 [15]),
      .O (\syn178132/FROM )
    );
    X_BUF \syn178132/YUSED (
      .I (\syn178132/GROM ),
      .O (syn178167)
    );
    X_BUF \syn178132/XUSED (
      .I (\syn178132/FROM ),
      .O (syn178132)
    );
    defparam C19488.INIT = 16'hFFEC;
    X_LUT4 C19488(
      .ADR0 (syn17067),
      .ADR1 (syn17118),
      .ADR2 (\bridge/conf_cache_line_size_out [0]),
      .ADR3 (syn17115),
      .O (\syn18717/GROM )
    );
    defparam C19537.INIT = 16'h8888;
    X_LUT4 C19537(
      .ADR0 (\bridge/conf_cache_line_size_out [4]),
      .ADR1 (syn17067),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn18717/FROM )
    );
    X_BUF \syn18717/YUSED (
      .I (\syn18717/GROM ),
      .O (syn178530)
    );
    X_BUF \syn18717/XUSED (
      .I (\syn18717/FROM ),
      .O (syn18717)
    );
    defparam C18864.INIT = 16'h4000;
    X_LUT4 C18864(
      .ADR0 (\bridge/in_reg_cbe_out [1]),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C294/N84/GROM )
    );
    defparam C18894.INIT = 16'h0080;
    X_LUT4 C18894(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/configuration/C1955 ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/in_reg_cbe_out [1]),
      .O (\bridge/configuration/C294/N84/FROM )
    );
    X_BUF \bridge/configuration/C294/N84/YUSED (
      .I (\bridge/configuration/C294/N84/GROM ),
      .O (\bridge/configuration/C299/N74 )
    );
    X_BUF \bridge/configuration/C294/N84/XUSED (
      .I (\bridge/configuration/C294/N84/FROM ),
      .O (\bridge/configuration/C294/N84 )
    );
    defparam C18856.INIT = 16'h0080;
    X_LUT4 C18856(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/configuration/C1989 ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/in_reg_cbe_out [2]),
      .O (\bridge/configuration/C294/N69/GROM )
    );
    defparam C18862.INIT = 16'h0080;
    X_LUT4 C18862(
      .ADR0 (\bridge/pciu_conf_offset_out [8]),
      .ADR1 (\bridge/configuration/C1955 ),
      .ADR2 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .ADR3 (\bridge/in_reg_cbe_out [2]),
      .O (\bridge/configuration/C294/N69/FROM )
    );
    X_BUF \bridge/configuration/C294/N69/YUSED (
      .I (\bridge/configuration/C294/N69/GROM ),
      .O (\bridge/configuration/C290/N54 )
    );
    X_BUF \bridge/configuration/C294/N69/XUSED (
      .I (\bridge/configuration/C294/N69/FROM ),
      .O (\bridge/configuration/C294/N69 )
    );
    defparam C18848.INIT = 16'h4000;
    X_LUT4 C18848(
      .ADR0 (\bridge/in_reg_cbe_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [8]),
      .ADR2 (\bridge/configuration/C1929 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C297/N69/GROM )
    );
    defparam C18851.INIT = 16'h2000;
    X_LUT4 C18851(
      .ADR0 (\bridge/configuration/C1951 ),
      .ADR1 (\bridge/in_reg_cbe_out [2]),
      .ADR2 (\bridge/pciu_conf_offset_out [8]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C297/N69/FROM )
    );
    X_BUF \bridge/configuration/C297/N69/YUSED (
      .I (\bridge/configuration/C297/N69/GROM ),
      .O (\bridge/configuration/C299/N29 )
    );
    X_BUF \bridge/configuration/C297/N69/XUSED (
      .I (\bridge/configuration/C297/N69/FROM ),
      .O (\bridge/configuration/C297/N69 )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_done_reg_clr/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_done_reg_clr/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_done_reg_clr_reg (
      .I (\bridge/pci_target_unit/del_sync/comp_done_reg_main ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_done_reg_clr/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_done_reg_clr )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_done_reg_clr/FFY/ASYNC_FF_GSR_OR_149 (
      .I0 (\bridge/pci_target_unit/del_sync/comp_done_reg_clr/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_done_reg_clr/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19825.INIT = 16'hF888;
    X_LUT4 C19825(
      .ADR0 (\bridge/configuration/C2308 ),
      .ADR1 (\bridge/configuration/wb_err_cs_bit31_24 [27]),
      .ADR2 (\bridge/configuration/C2302 ),
      .ADR3 (\bridge/configuration/wb_err_data [27]),
      .O (\syn177655/GROM )
    );
    defparam C19847.INIT = 16'hECA0;
    X_LUT4 C19847(
      .ADR0 (\bridge/configuration/wb_err_cs_bit31_24 [28]),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (\bridge/configuration/C2308 ),
      .ADR3 (\bridge/configuration/wb_err_data [28]),
      .O (\syn177655/FROM )
    );
    X_BUF \syn177655/YUSED (
      .I (\syn177655/GROM ),
      .O (syn177692)
    );
    X_BUF \syn177655/XUSED (
      .I (\syn177655/FROM ),
      .O (syn177655)
    );
    defparam C19809.INIT = 16'hECA0;
    X_LUT4 C19809(
      .ADR0 (syn17055),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [26]),
      .ADR2 (syn16928),
      .ADR3 (syn17745),
      .O (\syn177670/GROM )
    );
    defparam C19839.INIT = 16'hEAC0;
    X_LUT4 C19839(
      .ADR0 (syn17053),
      .ADR1 (syn17745),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [28]),
      .ADR3 (syn16928),
      .O (\syn177670/FROM )
    );
    X_BUF \syn177670/YUSED (
      .I (\syn177670/GROM ),
      .O (syn177749)
    );
    X_BUF \syn177670/XUSED (
      .I (\syn177670/FROM ),
      .O (syn177670)
    );
    defparam C19673.INIT = 16'hF888;
    X_LUT4 C19673(
      .ADR0 (\bridge/configuration/config_addr[16] ),
      .ADR1 (\bridge/configuration/C2296 ),
      .ADR2 (\bridge/configuration/wb_err_addr [16]),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn178058/GROM )
    );
    defparam C19686.INIT = 16'hF888;
    X_LUT4 C19686(
      .ADR0 (\bridge/configuration/wb_err_addr [17]),
      .ADR1 (\bridge/configuration/C2304 ),
      .ADR2 (\bridge/configuration/C2296 ),
      .ADR3 (\bridge/configuration/config_addr[17] ),
      .O (\syn178058/FROM )
    );
    X_BUF \syn178058/YUSED (
      .I (\syn178058/GROM ),
      .O (syn178096)
    );
    X_BUF \syn178058/XUSED (
      .I (\syn178058/FROM ),
      .O (syn178058)
    );
    defparam C19649.INIT = 16'hEAC0;
    X_LUT4 C19649(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [14]),
      .ADR2 (\bridge/configuration/C2318 ),
      .ADR3 (\bridge/configuration/pci_err_addr [14]),
      .O (\syn178131/GROM )
    );
    defparam C19664.INIT = 16'hF888;
    X_LUT4 C19664(
      .ADR0 (\bridge/configuration/C2318 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [15]),
      .ADR2 (\bridge/configuration/C2338 ),
      .ADR3 (\bridge/configuration/pci_err_addr [15]),
      .O (\syn178131/FROM )
    );
    X_BUF \syn178131/YUSED (
      .I (\syn178131/GROM ),
      .O (syn178166)
    );
    X_BUF \syn178131/XUSED (
      .I (\syn178131/FROM ),
      .O (syn178131)
    );
    defparam C19593.INIT = 16'hEAC0;
    X_LUT4 C19593(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [10]),
      .ADR1 (syn17074),
      .ADR2 (\bridge/configuration/wb_err_data [10]),
      .ADR3 (syn17745),
      .O (\syn18567/GROM )
    );
    defparam C19607.INIT = 16'hCC00;
    X_LUT4 C19607(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [11]),
      .ADR2 (VCC),
      .ADR3 (syn17745),
      .O (\syn18567/FROM )
    );
    X_BUF \syn18567/YUSED (
      .I (\syn18567/GROM ),
      .O (syn178293)
    );
    X_BUF \syn18567/XUSED (
      .I (\syn18567/FROM ),
      .O (syn18567)
    );
    defparam C19497.INIT = 16'hECA0;
    X_LUT4 C19497(
      .ADR0 (\bridge/configuration/wb_error_en ),
      .ADR1 (\bridge/configuration/wb_err_data [0]),
      .ADR2 (\bridge/configuration/C2308 ),
      .ADR3 (\bridge/configuration/C2302 ),
      .O (\syn177732/GROM )
    );
    defparam C19820.INIT = 16'hECA0;
    X_LUT4 C19820(
      .ADR0 (\bridge/configuration/wb_err_data [26]),
      .ADR1 (\bridge/configuration/C2308 ),
      .ADR2 (\bridge/configuration/C2302 ),
      .ADR3 (\bridge/configuration/wb_err_cs_bit31_24 [26]),
      .O (\syn177732/FROM )
    );
    X_BUF \syn177732/YUSED (
      .I (\syn177732/GROM ),
      .O (syn178515)
    );
    X_BUF \syn177732/XUSED (
      .I (\syn177732/FROM ),
      .O (syn177732)
    );
    defparam C19489.INIT = 16'hEAC0;
    X_LUT4 C19489(
      .ADR0 (\bridge/configuration/interrupt_line [0]),
      .ADR1 (syn17745),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [0]),
      .ADR3 (syn17083),
      .O (\syn18681/GROM )
    );
    defparam C19548.INIT = 16'hC0C0;
    X_LUT4 C19548(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [6]),
      .ADR2 (syn17745),
      .ADR3 (VCC),
      .O (\syn18681/FROM )
    );
    X_BUF \syn18681/YUSED (
      .I (\syn18681/GROM ),
      .O (syn178529)
    );
    X_BUF \syn18681/XUSED (
      .I (\syn18681/FROM ),
      .O (syn18681)
    );
    defparam C18929.INIT = 16'h7FFF;
    X_LUT4 C18929(
      .ADR0 (\CRT/ssvga_crtc/hcntr [0]),
      .ADR1 (\CRT/ssvga_crtc/hcntr [9]),
      .ADR2 (\CRT/ssvga_crtc/hcntr [7]),
      .ADR3 (\CRT/ssvga_crtc/hcntr [3]),
      .O (\syn20277/GROM )
    );
    defparam C18945.INIT = 16'h8001;
    X_LUT4 C18945(
      .ADR0 (\CRT/ssvga_crtc/hcntr [6]),
      .ADR1 (\CRT/ssvga_crtc/hcntr [3]),
      .ADR2 (\CRT/ssvga_crtc/hcntr [1]),
      .ADR3 (\CRT/ssvga_crtc/hcntr [4]),
      .O (\syn20277/FROM )
    );
    X_BUF \syn20277/YUSED (
      .I (\syn20277/GROM ),
      .O (syn179587)
    );
    X_BUF \syn20277/XUSED (
      .I (\syn20277/FROM ),
      .O (syn20277)
    );
    defparam C18865.INIT = 16'h4444;
    X_LUT4 C18865(
      .ADR0 (\bridge/in_reg_cbe_out [2]),
      .ADR1 (syn17097),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/configuration/C286/N54/GROM )
    );
    defparam C18914.INIT = 16'h2200;
    X_LUT4 C18914(
      .ADR0 (syn60110),
      .ADR1 (\bridge/in_reg_cbe_out [2]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C286/N54/FROM )
    );
    X_BUF \bridge/configuration/C286/N54/YUSED (
      .I (\bridge/configuration/C286/N54/GROM ),
      .O (\bridge/configuration/C285/N79 )
    );
    X_BUF \bridge/configuration/C286/N54/XUSED (
      .I (\bridge/configuration/C286/N54/FROM ),
      .O (\bridge/configuration/C286/N54 )
    );
    defparam C18785.INIT = 16'hFFFD;
    X_LUT4 C18785(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [0]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [2]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C262/GROM )
    );
    defparam C19482.INIT = 16'h0010;
    X_LUT4 C19482(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [0]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [2]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [1]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_sm/cur_state [3]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C262/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/C262/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C262/GROM ),
      .O (syn20490)
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/C262/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/C262/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C262 )
    );
    defparam C18697.INIT = 16'hF888;
    X_LUT4 C18697(
      .ADR0 (syn16983),
      .ADR1 (\bridge/configuration/pci_err_addr [5]),
      .ADR2 (syn16985),
      .ADR3 (\bridge/configuration/pci_err_data [5]),
      .O (\syn178394/GROM )
    );
    defparam C19541.INIT = 16'hEAC0;
    X_LUT4 C19541(
      .ADR0 (\bridge/conf_cache_line_size_out [5]),
      .ADR1 (\bridge/configuration/pci_err_data [5]),
      .ADR2 (syn17077),
      .ADR3 (syn17081),
      .O (\syn178394/FROM )
    );
    X_BUF \syn178394/YUSED (
      .I (\syn178394/GROM ),
      .O (syn180053)
    );
    X_BUF \syn178394/XUSED (
      .I (\syn178394/FROM ),
      .O (syn178394)
    );
    defparam C19842.INIT = 16'h8000;
    X_LUT4 C19842(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .O (\syn59929/GROM )
    );
    defparam C19916.INIT = 16'h3030;
    X_LUT4 C19916(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR3 (VCC),
      .O (\syn59929/FROM )
    );
    X_BUF \syn59929/YUSED (
      .I (\syn59929/GROM ),
      .O (syn177629)
    );
    X_BUF \syn59929/XUSED (
      .I (\syn59929/FROM ),
      .O (syn59929)
    );
    defparam C19578.INIT = 16'hEAC0;
    X_LUT4 C19578(
      .ADR0 (syn17077),
      .ADR1 (syn17081),
      .ADR2 (\bridge/conf_latency_tim_out [1]),
      .ADR3 (\bridge/configuration/pci_err_data [9]),
      .O (\syn178313/GROM )
    );
    X_BUF \syn178313/YUSED (
      .I (\syn178313/GROM ),
      .O (syn178313)
    );
    defparam C19498.INIT = 16'hECA0;
    X_LUT4 C19498(
      .ADR0 (\bridge/configuration/wb_img_ctrl1[0] ),
      .ADR1 (\bridge/configuration/C2292 ),
      .ADR2 (\bridge/configuration/C2326 ),
      .ADR3 (\bridge/configuration/int_prop_en ),
      .O (\syn178514/GROM )
    );
    X_BUF \syn178514/YUSED (
      .I (\syn178514/GROM ),
      .O (syn178514)
    );
    defparam C18954.INIT = 16'h0001;
    X_LUT4 C18954(
      .ADR0 (\CRT/ssvga_crtc/vcntr [1]),
      .ADR1 (\CRT/ssvga_crtc/vcntr [4]),
      .ADR2 (\CRT/ssvga_crtc/vcntr [3]),
      .ADR3 (\CRT/ssvga_crtc/vcntr [0]),
      .O (\syn179544/GROM )
    );
    X_BUF \syn179544/YUSED (
      .I (\syn179544/GROM ),
      .O (syn179544)
    );
    defparam C18778.INIT = 16'h0302;
    X_LUT4 C18778(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/norm_access_to_conf_reg ),
      .ADR1 (\bridge/out_bckp_devsel_out ),
      .ADR2 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/cnf_progress ),
      .O (\syn19914/GROM )
    );
    defparam C19149.INIT = 16'hEECC;
    X_LUT4 C19149(
      .ADR0 (\bridge/pci_target_unit/pci_target_sm/wr_progress ),
      .ADR1 (\bridge/pci_target_unit/pci_target_sm/cnf_progress ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pcit_sm_bc0_out ),
      .O (\syn19914/FROM )
    );
    X_BUF \syn19914/YUSED (
      .I (\syn19914/GROM ),
      .O (syn17106)
    );
    X_BUF \syn19914/XUSED (
      .I (\syn19914/FROM ),
      .O (syn19914)
    );
    defparam C19587.INIT = 16'h8080;
    X_LUT4 C19587(
      .ADR0 (\bridge/configuration/pci_error_rty_exp_set ),
      .ADR1 (\bridge/configuration/C2340 ),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR3 (VCC),
      .O (\syn17080/GROM )
    );
    defparam C19595.INIT = 16'hA0A0;
    X_LUT4 C19595(
      .ADR0 (\bridge/configuration/C2308 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C92 ),
      .ADR3 (VCC),
      .O (\syn17080/FROM )
    );
    X_BUF \syn17080/YUSED (
      .I (\syn17080/GROM ),
      .O (syn18585)
    );
    X_BUF \syn17080/XUSED (
      .I (\syn17080/FROM ),
      .O (syn17080)
    );
    defparam C18955.INIT = 16'hFFFE;
    X_LUT4 C18955(
      .ADR0 (\CRT/ssvga_crtc/vcntr [6]),
      .ADR1 (\CRT/ssvga_crtc/vcntr [7]),
      .ADR2 (\CRT/ssvga_crtc/vcntr [8]),
      .ADR3 (\CRT/ssvga_crtc/vcntr [5]),
      .O (\syn16988/GROM )
    );
    X_BUF \syn16988/YUSED (
      .I (\syn16988/GROM ),
      .O (syn16988)
    );
    defparam C18947.INIT = 16'h0AAA;
    X_LUT4 C18947(
      .ADR0 (syn16982),
      .ADR1 (VCC),
      .ADR2 (syn16991),
      .ADR3 (syn16988),
      .O (\N12163/GROM )
    );
    defparam C18952.INIT = 16'h4040;
    X_LUT4 C18952(
      .ADR0 (syn16988),
      .ADR1 (syn179544),
      .ADR2 (syn179548),
      .ADR3 (VCC),
      .O (\N12163/FROM )
    );
    X_BUF \N12163/YUSED (
      .I (\N12163/GROM ),
      .O (N12162)
    );
    X_BUF \N12163/XUSED (
      .I (\N12163/FROM ),
      .O (N12163)
    );
    defparam C18939.INIT = 16'h5050;
    X_LUT4 C18939(
      .ADR0 (\CRT/ssvga_crtc/line_end2 ),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/line_end1 ),
      .ADR3 (VCC),
      .O (\N12152/GROM )
    );
    X_BUF \N12152/YUSED (
      .I (\N12152/GROM ),
      .O (N12152)
    );
    defparam C18891.INIT = 16'hFFAF;
    X_LUT4 C18891(
      .ADR0 (\bridge/pciu_conf_offset_out [4]),
      .ADR1 (VCC),
      .ADR2 (\bridge/pciu_conf_offset_out [3]),
      .ADR3 (\bridge/pciu_conf_offset_out [7]),
      .O (\syn20367/GROM )
    );
    defparam C18893.INIT = 16'h00A7;
    X_LUT4 C18893(
      .ADR0 (\bridge/pciu_conf_offset_out [7]),
      .ADR1 (\bridge/pciu_conf_offset_out [4]),
      .ADR2 (\bridge/pciu_conf_offset_out [6]),
      .ADR3 (\bridge/pciu_conf_offset_out [5]),
      .O (\syn20367/FROM )
    );
    X_BUF \syn20367/YUSED (
      .I (\syn20367/GROM ),
      .O (syn20368)
    );
    X_BUF \syn20367/XUSED (
      .I (\syn20367/FROM ),
      .O (syn20367)
    );
    defparam C17899.INIT = 16'h5410;
    X_LUT4 C17899(
      .ADR0 (syn19562),
      .ADR1 (syn19555),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C960 ),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .O (\N12312/GROM )
    );
    defparam C18838.INIT = 16'h4000;
    X_LUT4 C18838(
      .ADR0 (syn19562),
      .ADR1 (\bridge/configuration/pci_error_en ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C981 ),
      .ADR3 (syn19555),
      .O (\N12312/FROM )
    );
    X_BUF \N12312/YUSED (
      .I (\N12312/GROM ),
      .O (syn182107)
    );
    X_BUF \N12312/XUSED (
      .I (\N12312/FROM ),
      .O (N12312)
    );
    defparam C19836.INIT = 16'h8888;
    X_LUT4 C19836(
      .ADR0 (\bridge/conf_pci_ba1_out [15]),
      .ADR1 (\bridge/conf_pci_am1_out [15]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn17054/GROM )
    );
    X_BUF \syn17054/YUSED (
      .I (\syn17054/GROM ),
      .O (syn17054)
    );
    defparam C19748.INIT = 16'hECA0;
    X_LUT4 C19748(
      .ADR0 (syn16928),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [22]),
      .ADR2 (syn17059),
      .ADR3 (syn17745),
      .O (\syn177790/GROM )
    );
    defparam C19804.INIT = 16'hEAC0;
    X_LUT4 C19804(
      .ADR0 (syn17056),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [25]),
      .ADR2 (syn17745),
      .ADR3 (syn16928),
      .O (\syn177790/FROM )
    );
    X_BUF \syn177790/YUSED (
      .I (\syn177790/GROM ),
      .O (syn177902)
    );
    X_BUF \syn177790/XUSED (
      .I (\syn177790/FROM ),
      .O (syn177790)
    );
    defparam C18796.INIT = 16'hF888;
    X_LUT4 C18796(
      .ADR0 (syn60110),
      .ADR1 (\bridge/conf_pci_mem_io1_out ),
      .ADR2 (\bridge/configuration/pci_error_en ),
      .ADR3 (\bridge/configuration/C1973 ),
      .O (\bridge/configuration/C286/N99/GROM )
    );
    defparam C18907.INIT = 16'h0A00;
    X_LUT4 C18907(
      .ADR0 (syn60110),
      .ADR1 (VCC),
      .ADR2 (\bridge/in_reg_cbe_out [1]),
      .ADR3 (\bridge/pci_target_unit/pci_target_sm/S_345/cell0 ),
      .O (\bridge/configuration/C286/N99/FROM )
    );
    X_BUF \bridge/configuration/C286/N99/YUSED (
      .I (\bridge/configuration/C286/N99/GROM ),
      .O (syn179851)
    );
    X_BUF \bridge/configuration/C286/N99/XUSED (
      .I (\bridge/configuration/C286/N99/FROM ),
      .O (\bridge/configuration/C286/N99 )
    );
    defparam C19861.INIT = 16'hE0A0;
    X_LUT4 C19861(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/conf_wb_ba1_out [17]),
      .ADR2 (\bridge/conf_wb_am1_out [17]),
      .ADR3 (\bridge/configuration/C2322 ),
      .O (\syn17856/GROM )
    );
    defparam C19878.INIT = 16'hE0C0;
    X_LUT4 C19878(
      .ADR0 (\bridge/configuration/C2322 ),
      .ADR1 (\bridge/configuration/C2320 ),
      .ADR2 (\bridge/conf_wb_am1_out [18]),
      .ADR3 (\bridge/conf_wb_ba1_out [18]),
      .O (\syn17856/FROM )
    );
    X_BUF \syn17856/YUSED (
      .I (\syn17856/GROM ),
      .O (syn17894)
    );
    X_BUF \syn17856/XUSED (
      .I (\syn17856/FROM ),
      .O (syn17856)
    );
    defparam C19781.INIT = 16'hF888;
    X_LUT4 C19781(
      .ADR0 (\bridge/configuration/pci_err_addr [24]),
      .ADR1 (\bridge/configuration/C2338 ),
      .ADR2 (\bridge/configuration/C2370 ),
      .ADR3 (\bridge/conf_pci_ba0_out [12]),
      .O (\syn177693/GROM )
    );
    defparam C19826.INIT = 16'hF888;
    X_LUT4 C19826(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/pci_err_addr [27]),
      .ADR2 (\bridge/conf_pci_ba0_out [15]),
      .ADR3 (\bridge/configuration/C2370 ),
      .O (\syn177693/FROM )
    );
    X_BUF \syn177693/YUSED (
      .I (\syn177693/GROM ),
      .O (syn177815)
    );
    X_BUF \syn177693/XUSED (
      .I (\syn177693/FROM ),
      .O (syn177693)
    );
    defparam C19757.INIT = 16'hEAC0;
    X_LUT4 C19757(
      .ADR0 (\bridge/configuration/pci_base_addr0 [22]),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [22]),
      .ADR2 (\bridge/configuration/C2320 ),
      .ADR3 (\bridge/configuration/C2370 ),
      .O (\syn177857/GROM )
    );
    defparam C19772.INIT = 16'hEAC0;
    X_LUT4 C19772(
      .ADR0 (\bridge/configuration/pci_base_addr0 [23]),
      .ADR1 (\bridge/configuration/wb_addr_mask1 [23]),
      .ADR2 (\bridge/configuration/C2320 ),
      .ADR3 (\bridge/configuration/C2370 ),
      .O (\syn177857/FROM )
    );
    X_BUF \syn177857/YUSED (
      .I (\syn177857/GROM ),
      .O (syn177890)
    );
    X_BUF \syn177857/XUSED (
      .I (\syn177857/FROM ),
      .O (syn177857)
    );
    defparam C19934.INIT = 16'hC000;
    X_LUT4 C19934(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR2 (syn177397),
      .ADR3 (syn177396),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C116/GROM )
    );
    X_BUF \bridge/wishbone_slave_unit/wb_addr_dec/C0/C116/YUSED (
      .I (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C116/GROM ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C116 )
    );
    defparam C19862.INIT = 16'hEAC0;
    X_LUT4 C19862(
      .ADR0 (\bridge/conf_pci_am1_out [17]),
      .ADR1 (\bridge/configuration/C2354 ),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [29]),
      .ADR3 (\bridge/configuration/C2356 ),
      .O (\syn177574/GROM )
    );
    defparam C19872.INIT = 16'hEAC0;
    X_LUT4 C19872(
      .ADR0 (\bridge/conf_pci_am1_out [18]),
      .ADR1 (\bridge/configuration/C2354 ),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [30]),
      .ADR3 (\bridge/configuration/C2356 ),
      .O (\syn177574/FROM )
    );
    X_BUF \syn177574/YUSED (
      .I (\syn177574/GROM ),
      .O (syn177614)
    );
    X_BUF \syn177574/XUSED (
      .I (\syn177574/FROM ),
      .O (syn177574)
    );
    defparam C19782.INIT = 16'hA8A0;
    X_LUT4 C19782(
      .ADR0 (\bridge/conf_wb_am1_out [12]),
      .ADR1 (\bridge/conf_wb_ba1_out [12]),
      .ADR2 (\bridge/configuration/C2320 ),
      .ADR3 (\bridge/configuration/C2322 ),
      .O (\syn18010/GROM )
    );
    defparam C19813.INIT = 16'hE0C0;
    X_LUT4 C19813(
      .ADR0 (\bridge/configuration/C2322 ),
      .ADR1 (\bridge/configuration/C2320 ),
      .ADR2 (\bridge/conf_wb_am1_out [14]),
      .ADR3 (\bridge/conf_wb_ba1_out [14]),
      .O (\syn18010/FROM )
    );
    X_BUF \syn18010/YUSED (
      .I (\syn18010/GROM ),
      .O (syn18086)
    );
    X_BUF \syn18010/XUSED (
      .I (\syn18010/FROM ),
      .O (syn18010)
    );
    defparam C19758.INIT = 16'hEAC0;
    X_LUT4 C19758(
      .ADR0 (\bridge/configuration/C2338 ),
      .ADR1 (\bridge/configuration/wb_tran_addr1 [22]),
      .ADR2 (\bridge/configuration/C2318 ),
      .ADR3 (\bridge/configuration/pci_err_addr [22]),
      .O (\syn177856/GROM )
    );
    defparam C19773.INIT = 16'hEAC0;
    X_LUT4 C19773(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [23]),
      .ADR1 (\bridge/configuration/C2338 ),
      .ADR2 (\bridge/configuration/pci_err_addr [23]),
      .ADR3 (\bridge/configuration/C2318 ),
      .O (\syn177856/FROM )
    );
    X_BUF \syn177856/YUSED (
      .I (\syn177856/GROM ),
      .O (syn177889)
    );
    X_BUF \syn177856/XUSED (
      .I (\syn177856/FROM ),
      .O (syn177856)
    );
    defparam C19919.INIT = 16'h8000;
    X_LUT4 C19919(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR3 (syn177475),
      .O (\syn60060/GROM )
    );
    defparam C19954.INIT = 16'h5500;
    X_LUT4 C19954(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .O (\syn60060/FROM )
    );
    X_BUF \syn60060/YUSED (
      .I (\syn60060/GROM ),
      .O (syn177458)
    );
    X_BUF \syn60060/XUSED (
      .I (\syn60060/FROM ),
      .O (syn60060)
    );
    defparam C19855.INIT = 16'hAA00;
    X_LUT4 C19855(
      .ADR0 (syn16930),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_pci_ba0_out [17]),
      .O (\syn177609/GROM )
    );
    defparam C19860.INIT = 16'hEAC0;
    X_LUT4 C19860(
      .ADR0 (\bridge/conf_pci_ba0_out [17]),
      .ADR1 (\bridge/configuration/C2338 ),
      .ADR2 (\bridge/configuration/pci_err_addr [29]),
      .ADR3 (\bridge/configuration/C2370 ),
      .O (\syn177609/FROM )
    );
    X_BUF \syn177609/YUSED (
      .I (\syn177609/GROM ),
      .O (syn17912)
    );
    X_BUF \syn177609/XUSED (
      .I (\syn177609/FROM ),
      .O (syn177609)
    );
    defparam C19679.INIT = 16'hECA0;
    X_LUT4 C19679(
      .ADR0 (\bridge/configuration/C2318 ),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (\bridge/configuration/wb_tran_addr1 [16]),
      .ADR3 (\bridge/configuration/wb_err_data [16]),
      .O (\syn178055/GROM )
    );
    defparam C19692.INIT = 16'hEAC0;
    X_LUT4 C19692(
      .ADR0 (\bridge/configuration/C2318 ),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (\bridge/configuration/wb_err_data [17]),
      .ADR3 (\bridge/configuration/wb_tran_addr1 [17]),
      .O (\syn178055/FROM )
    );
    X_BUF \syn178055/YUSED (
      .I (\syn178055/GROM ),
      .O (syn178093)
    );
    X_BUF \syn178055/XUSED (
      .I (\syn178055/FROM ),
      .O (syn178055)
    );
    defparam C18959.INIT = 16'hFF7F;
    X_LUT4 C18959(
      .ADR0 (\CRT/ssvga_crtc/hcntr [2]),
      .ADR1 (\CRT/ssvga_crtc/hcntr [6]),
      .ADR2 (\CRT/ssvga_crtc/hcntr [5]),
      .ADR3 (\CRT/ssvga_crtc/hcntr [8]),
      .O (\syn48756/GROM )
    );
    X_BUF \syn48756/YUSED (
      .I (\syn48756/GROM ),
      .O (syn48756)
    );
    defparam C19960.INIT = 16'h5500;
    X_LUT4 C19960(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .O (\syn50321/GROM )
    );
    X_BUF \syn50321/YUSED (
      .I (\syn50321/GROM ),
      .O (syn50321)
    );
    defparam C19848.INIT = 16'hECCC;
    X_LUT4 C19848(
      .ADR0 (\bridge/conf_wb_ba1_out [16]),
      .ADR1 (\bridge/configuration/C2368 ),
      .ADR2 (\bridge/configuration/C2322 ),
      .ADR3 (\bridge/conf_wb_am1_out [16]),
      .O (\syn177657/GROM )
    );
    defparam C19851.INIT = 16'hF888;
    X_LUT4 C19851(
      .ADR0 (\bridge/configuration/C2320 ),
      .ADR1 (\bridge/conf_wb_am1_out [16]),
      .ADR2 (\bridge/conf_pci_ba0_out [16]),
      .ADR3 (\bridge/configuration/C2370 ),
      .O (\syn177657/FROM )
    );
    X_BUF \syn177657/YUSED (
      .I (\syn177657/GROM ),
      .O (syn177654)
    );
    X_BUF \syn177657/XUSED (
      .I (\syn177657/FROM ),
      .O (syn177657)
    );
    defparam C19784.INIT = 16'hF888;
    X_LUT4 C19784(
      .ADR0 (\bridge/configuration/pci_err_cs_bit31_24 [24]),
      .ADR1 (\bridge/configuration/C2340 ),
      .ADR2 (\bridge/configuration/pci_err_data [24]),
      .ADR3 (\bridge/configuration/C2334 ),
      .O (\syn177778/GROM )
    );
    defparam C19794.INIT = 16'hECA0;
    X_LUT4 C19794(
      .ADR0 (\bridge/configuration/pci_err_data [25]),
      .ADR1 (\bridge/configuration/C2340 ),
      .ADR2 (\bridge/configuration/C2334 ),
      .ADR3 (\bridge/configuration/pci_err_cs_bit31_24 [25]),
      .O (\syn177778/FROM )
    );
    X_BUF \syn177778/YUSED (
      .I (\syn177778/GROM ),
      .O (syn177819)
    );
    X_BUF \syn177778/XUSED (
      .I (\syn177778/FROM ),
      .O (syn177778)
    );
    defparam C19776.INIT = 16'hA0A0;
    X_LUT4 C19776(
      .ADR0 (syn16930),
      .ADR1 (VCC),
      .ADR2 (\bridge/conf_pci_ba0_out [12]),
      .ADR3 (VCC),
      .O (\syn17990/GROM )
    );
    defparam C19827.INIT = 16'hC0C0;
    X_LUT4 C19827(
      .ADR0 (VCC),
      .ADR1 (syn16930),
      .ADR2 (\bridge/conf_pci_ba0_out [15]),
      .ADR3 (VCC),
      .O (\syn17990/FROM )
    );
    X_BUF \syn17990/YUSED (
      .I (\syn17990/GROM ),
      .O (syn18104)
    );
    X_BUF \syn17990/XUSED (
      .I (\syn17990/FROM ),
      .O (syn17990)
    );
    defparam C18888.INIT = 16'hF7F4;
    X_LUT4 C18888(
      .ADR0 (\bridge/pciu_conf_offset_out [6]),
      .ADR1 (\bridge/pciu_conf_offset_out [4]),
      .ADR2 (\bridge/pciu_conf_offset_out [3]),
      .ADR3 (\bridge/pciu_conf_offset_out [5]),
      .O (\syn60089/GROM )
    );
    defparam C18916.INIT = 16'h0020;
    X_LUT4 C18916(
      .ADR0 (\bridge/pciu_conf_offset_out [2]),
      .ADR1 (\bridge/pciu_conf_offset_out [3]),
      .ADR2 (\bridge/pciu_conf_offset_out [4]),
      .ADR3 (\bridge/pciu_conf_offset_out [5]),
      .O (\syn60089/FROM )
    );
    X_BUF \syn60089/YUSED (
      .I (\syn60089/GROM ),
      .O (syn20360)
    );
    X_BUF \syn60089/XUSED (
      .I (\syn60089/FROM ),
      .O (syn60089)
    );
    defparam C19945.INIT = 16'h84CC;
    X_LUT4 C19945(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [26]),
      .ADR1 (syn60046),
      .ADR2 (\bridge/conf_wb_ba1_out [14]),
      .ADR3 (\bridge/conf_wb_am1_out [14]),
      .O (\syn60045/GROM )
    );
    defparam C19966.INIT = 16'hBB77;
    X_LUT4 C19966(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [26]),
      .ADR1 (\bridge/conf_wb_am1_out [14]),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_wb_ba1_out [14]),
      .O (\syn60045/FROM )
    );
    X_BUF \syn60045/YUSED (
      .I (\syn60045/GROM ),
      .O (syn177393)
    );
    X_BUF \syn60045/XUSED (
      .I (\syn60045/FROM ),
      .O (syn60045)
    );
    defparam C19881.INIT = 16'hEAC0;
    X_LUT4 C19881(
      .ADR0 (\bridge/configuration/C2308 ),
      .ADR1 (\bridge/configuration/C2302 ),
      .ADR2 (\bridge/configuration/wb_err_data [30]),
      .ADR3 (\bridge/configuration/wb_err_cs_bit31_24 [30]),
      .O (\syn177568/GROM )
    );
    X_BUF \syn177568/YUSED (
      .I (\syn177568/GROM ),
      .O (syn177568)
    );
    defparam C19857.INIT = 16'hECA0;
    X_LUT4 C19857(
      .ADR0 (syn17745),
      .ADR1 (\bridge/configuration/status_bit15_11 [13]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [29]),
      .ADR3 (syn24559),
      .O (\syn177585/GROM )
    );
    defparam C19871.INIT = 16'hEAC0;
    X_LUT4 C19871(
      .ADR0 (\bridge/configuration/status_bit15_11 [14]),
      .ADR1 (syn17745),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbr_data_out [30]),
      .ADR3 (syn24559),
      .O (\syn177585/FROM )
    );
    X_BUF \syn177585/YUSED (
      .I (\syn177585/GROM ),
      .O (syn177624)
    );
    X_BUF \syn177585/XUSED (
      .I (\syn177585/FROM ),
      .O (syn177585)
    );
    defparam C19793.INIT = 16'hEAC0;
    X_LUT4 C19793(
      .ADR0 (\bridge/configuration/pci_tran_addr1 [25]),
      .ADR1 (\bridge/configuration/C2356 ),
      .ADR2 (\bridge/conf_pci_am1_out [13]),
      .ADR3 (\bridge/configuration/C2354 ),
      .O (\syn177738/GROM )
    );
    defparam C19814.INIT = 16'hF888;
    X_LUT4 C19814(
      .ADR0 (\bridge/conf_pci_am1_out [14]),
      .ADR1 (\bridge/configuration/C2356 ),
      .ADR2 (\bridge/configuration/pci_tran_addr1 [26]),
      .ADR3 (\bridge/configuration/C2354 ),
      .O (\syn177738/FROM )
    );
    X_BUF \syn177738/YUSED (
      .I (\syn177738/GROM ),
      .O (syn177779)
    );
    X_BUF \syn177738/XUSED (
      .I (\syn177738/FROM ),
      .O (syn177738)
    );
    defparam C19777.INIT = 16'hF000;
    X_LUT4 C19777(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/conf_pci_ba1_out [12]),
      .ADR3 (\bridge/conf_pci_am1_out [12]),
      .O (\syn17057/GROM )
    );
    X_BUF \syn17057/YUSED (
      .I (\syn17057/GROM ),
      .O (syn17057)
    );
    defparam C18993.INIT = 16'hDDDD;
    X_LUT4 C18993(
      .ADR0 (N_LED),
      .ADR1 (\CRT/fifo_wr_en ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\N12065/GROM )
    );
    defparam C19054.INIT = 16'hFFCC;
    X_LUT4 C19054(
      .ADR0 (VCC),
      .ADR1 (\CRT/fifo_wr_en ),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_wbm_if/frame_read ),
      .O (\N12065/FROM )
    );
    X_BUF \N12065/YUSED (
      .I (\N12065/GROM ),
      .O (N12092)
    );
    X_BUF \N12065/XUSED (
      .I (\N12065/FROM ),
      .O (N12065)
    );
    defparam C18897.INIT = 16'hAA00;
    X_LUT4 C18897(
      .ADR0 (\bridge/pciu_conf_offset_out [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pciu_conf_offset_out [6]),
      .O (\syn17004/GROM )
    );
    defparam C18901.INIT = 16'h00CC;
    X_LUT4 C18901(
      .ADR0 (VCC),
      .ADR1 (\bridge/pciu_conf_offset_out [7]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pciu_conf_offset_out [6]),
      .O (\syn17004/FROM )
    );
    X_BUF \syn17004/YUSED (
      .I (\syn17004/GROM ),
      .O (syn17043)
    );
    X_BUF \syn17004/XUSED (
      .I (\syn17004/FROM ),
      .O (syn17004)
    );
    defparam C19875.INIT = 16'h0800;
    X_LUT4 C19875(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .O (\syn177501/GROM )
    );
    defparam C19931.INIT = 16'h0C00;
    X_LUT4 C19931(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .O (\syn177501/FROM )
    );
    X_BUF \syn177501/YUSED (
      .I (\syn177501/GROM ),
      .O (syn177548)
    );
    X_BUF \syn177501/XUSED (
      .I (\syn177501/FROM ),
      .O (syn177501)
    );
    defparam C19787.INIT = 16'hF888;
    X_LUT4 C19787(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [24]),
      .ADR1 (\bridge/configuration/C2318 ),
      .ADR2 (\bridge/configuration/wb_err_cs_bit31_24 [24]),
      .ADR3 (\bridge/configuration/C2308 ),
      .O (\syn177608/GROM )
    );
    defparam C19866.INIT = 16'hECA0;
    X_LUT4 C19866(
      .ADR0 (\bridge/configuration/C2308 ),
      .ADR1 (\bridge/configuration/C2318 ),
      .ADR2 (\bridge/configuration/wb_err_cs_bit31_24 [29]),
      .ADR3 (\bridge/configuration/wb_tran_addr1 [29]),
      .O (\syn177608/FROM )
    );
    X_BUF \syn177608/YUSED (
      .I (\syn177608/GROM ),
      .O (syn177814)
    );
    X_BUF \syn177608/XUSED (
      .I (\syn177608/FROM ),
      .O (syn177608)
    );
    defparam C19877.INIT = 16'hECA0;
    X_LUT4 C19877(
      .ADR0 (\bridge/conf_pci_ba0_out [18]),
      .ADR1 (\bridge/configuration/pci_err_addr [30]),
      .ADR2 (\bridge/configuration/C2370 ),
      .ADR3 (\bridge/configuration/C2338 ),
      .O (\syn177569/GROM )
    );
    X_BUF \syn177569/YUSED (
      .I (\syn177569/GROM ),
      .O (syn177569)
    );
    defparam C19797.INIT = 16'hF888;
    X_LUT4 C19797(
      .ADR0 (\bridge/configuration/pci_err_addr [25]),
      .ADR1 (\bridge/configuration/C2338 ),
      .ADR2 (\bridge/configuration/wb_err_cs_bit31_24 [25]),
      .ADR3 (\bridge/configuration/C2308 ),
      .O (\syn177656/GROM )
    );
    defparam C19852.INIT = 16'hF888;
    X_LUT4 C19852(
      .ADR0 (\bridge/configuration/wb_tran_addr1 [28]),
      .ADR1 (\bridge/configuration/C2318 ),
      .ADR2 (\bridge/configuration/C2338 ),
      .ADR3 (\bridge/configuration/pci_err_addr [28]),
      .O (\syn177656/FROM )
    );
    X_BUF \syn177656/YUSED (
      .I (\syn177656/GROM ),
      .O (syn177772)
    );
    X_BUF \syn177656/XUSED (
      .I (\syn177656/FROM ),
      .O (syn177656)
    );
    defparam C19798.INIT = 16'hECEC;
    X_LUT4 C19798(
      .ADR0 (\bridge/configuration/C2302 ),
      .ADR1 (\bridge/configuration/C2368 ),
      .ADR2 (\bridge/configuration/wb_err_data [25]),
      .ADR3 (VCC),
      .O (\syn17115/GROM )
    );
    defparam C19808.INIT = 16'h8888;
    X_LUT4 C19808(
      .ADR0 (syn177631),
      .ADR1 (\bridge/configuration/C2368 ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn17115/FROM )
    );
    X_BUF \syn17115/YUSED (
      .I (\syn17115/GROM ),
      .O (syn177771)
    );
    X_BUF \syn17115/XUSED (
      .I (\syn17115/FROM ),
      .O (syn17115)
    );
    X_INV \bridge/configuration/wb_error_en/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/wb_error_en/SRNOT )
    );
    X_FF \bridge/configuration/wb_err_cs_bit0_reg (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C298/N3 ),
      .SET (GND),
      .RST (\bridge/configuration/wb_error_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/wb_error_en )
    );
    X_OR2 \bridge/configuration/wb_error_en/FFY/ASYNC_FF_GSR_OR_150 (
      .I0 (\bridge/configuration/wb_error_en/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/wb_error_en/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C19991.INIT = 16'hB7DE;
    X_LUT4 C19991(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr_plus1 [6]),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [7]),
      .ADR2 (\CRT/ssvga_fifo/gray_read_ptr [8]),
      .ADR3 (\CRT/ssvga_fifo/gray_read_ptr [9]),
      .O (\syn177260/GROM )
    );
    defparam C20012.INIT = 16'h0C03;
    X_LUT4 C20012(
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr [7]),
      .ADR2 (\CRT/ssvga_fifo/gray_read_ptr [0]),
      .ADR3 (\CRT/ssvga_fifo/gray_read_ptr [9]),
      .O (\syn177260/FROM )
    );
    X_BUF \syn177260/YUSED (
      .I (\syn177260/GROM ),
      .O (syn177317)
    );
    X_BUF \syn177260/XUSED (
      .I (\syn177260/FROM ),
      .O (syn177260)
    );
    defparam C19959.INIT = 16'hF000;
    X_LUT4 C19959(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .O (\syn177541/GROM )
    );
    X_BUF \syn177541/YUSED (
      .I (\syn177541/GROM ),
      .O (syn177541)
    );
    defparam C19799.INIT = 16'hF000;
    X_LUT4 C19799(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/configuration/wb_err_addr [25]),
      .ADR3 (\bridge/configuration/C2304 ),
      .O (\syn18051/GROM )
    );
    X_BUF \syn18051/YUSED (
      .I (\syn18051/GROM ),
      .O (syn18051)
    );
    defparam C18999.INIT = 16'hAAFF;
    X_LUT4 C18999(
      .ADR0 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ssvga_en ),
      .O (\CRT/ssvga_fifo/C6/N6/GROM )
    );
    defparam C20000.INIT = 16'hDD88;
    X_LUT4 C20000(
      .ADR0 (\CRT/ssvga_fifo/S_45/cell0 ),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [0]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr [0]),
      .O (\CRT/ssvga_fifo/C6/N6/FROM )
    );
    X_BUF \CRT/ssvga_fifo/C6/N6/YUSED (
      .I (\CRT/ssvga_fifo/C6/N6/GROM ),
      .O (N12082)
    );
    X_BUF \CRT/ssvga_fifo/C6/N6/XUSED (
      .I (\CRT/ssvga_fifo/C6/N6/FROM ),
      .O (\CRT/ssvga_fifo/C6/N6 )
    );
    defparam C19992.INIT = 16'h9966;
    X_LUT4 C19992(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr_plus1 [4]),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [5]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/gray_read_ptr [6]),
      .O (\syn176894/GROM )
    );
    defparam C19993.INIT = 16'h9966;
    X_LUT4 C19993(
      .ADR0 (\CRT/ssvga_fifo/wr_ptr_plus1 [6]),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [5]),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/gray_read_ptr [7]),
      .O (\syn176894/FROM )
    );
    X_BUF \syn176894/YUSED (
      .I (\syn176894/GROM ),
      .O (syn176895)
    );
    X_BUF \syn176894/XUSED (
      .I (\syn176894/FROM ),
      .O (syn176894)
    );
    defparam C19976.INIT = 16'h0C00;
    X_LUT4 C19976(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [1]),
      .ADR2 (syn177324),
      .ADR3 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [2]),
      .O (\syn177406/GROM )
    );
    defparam C19982.INIT = 16'h8888;
    X_LUT4 C19982(
      .ADR0 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [0]),
      .ADR1 (\bridge/wishbone_slave_unit/wishbone_slave/c_state [1]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\syn177406/FROM )
    );
    X_BUF \syn177406/YUSED (
      .I (\syn177406/GROM ),
      .O (syn17686)
    );
    X_BUF \syn177406/XUSED (
      .I (\syn177406/FROM ),
      .O (syn177406)
    );
    defparam C19888.INIT = 16'hCE00;
    X_LUT4 C19888(
      .ADR0 (syn177440),
      .ADR1 (\bridge/configuration/C2368 ),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR3 (syn24500),
      .O (\syn177563/GROM )
    );
    defparam C19956.INIT = 16'h0505;
    X_LUT4 C19956(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .ADR3 (VCC),
      .O (\syn177563/FROM )
    );
    X_BUF \syn177563/YUSED (
      .I (\syn177563/GROM ),
      .O (syn48759)
    );
    X_BUF \syn177563/XUSED (
      .I (\syn177563/FROM ),
      .O (syn177563)
    );
    defparam C19897.INIT = 16'h5FFF;
    X_LUT4 C19897(
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR1 (VCC),
      .ADR2 (syn177396),
      .ADR3 (syn177397),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C112/GROM )
    );
    defparam C19928.INIT = 16'hA000;
    X_LUT4 C19928(
      .ADR0 (syn177397),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR3 (syn177396),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C112/FROM )
    );
    X_BUF \bridge/wishbone_slave_unit/wb_addr_dec/C0/C112/YUSED (
      .I (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C112/GROM ),
      .O (syn59978)
    );
    X_BUF \bridge/wishbone_slave_unit/wb_addr_dec/C0/C112/XUSED (
      .I (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C112/FROM ),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/C0/C112 )
    );
    defparam \bridge/parity_checker/par_gen/C72 .INIT = 16'hF0AA;
    X_LUT4 \bridge/parity_checker/par_gen/C72 (
      .ADR0 (\bridge/parity_checker/par_gen/syn143 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/parity_checker/par_out_only ),
      .ADR3 (\bridge/out_bckp_cbe_en_out ),
      .O (\bridge/pci_mux_par_in/GROM )
    );
    X_BUF \bridge/pci_mux_par_in/YUSED (
      .I (\bridge/pci_mux_par_in/GROM ),
      .O (\bridge/pci_mux_par_in )
    );
    X_INV \bridge/configuration/pci_base_addr0<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr0[21]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N79 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [20])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N79 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [21])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr0<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr0[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [12])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [13])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync/sync_req_comp_pending/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/sync_req_comp_pending/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_sync/sync_data_out_reg<0> (
      .I (\bridge/pciu_pci_drcomp_pending_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/sync_req_comp_pending/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/sync_req_comp_pending )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/sync_req_comp_pending/FFY/ASYNC_FF_GSR_OR_151 (
      .I0 (\bridge/pci_target_unit/del_sync/sync_req_comp_pending/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/sync_req_comp_pending/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_sync/sync_data_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_comp_pending_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending/FFY/ASYNC_FF_GSR_OR_152 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/sync_req_comp_pending/FFY/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/conf_pci_ba0_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_ba0_out[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<30> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N34 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba0_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba0_out [18])
    );
    X_OR2 \bridge/conf_pci_ba0_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba0_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba0_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<31> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N34 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba0_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba0_out [19])
    );
    X_OR2 \bridge/conf_pci_ba0_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba0_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba0_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr0<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr0[23]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N79 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [22])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N79 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [23])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr0<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr0[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [14])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N99 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [15])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_ONE \bridge/conf_wb_err_pending_out/LOGIC_ONE_153 (
      .O (\bridge/conf_wb_err_pending_out/LOGIC_ONE )
    );
    X_FF \bridge/configuration/wb_err_cs_bit10_8_reg3<8> (
      .I (\bridge/conf_wb_err_pending_out/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12237),
      .SET (GND),
      .RST (\bridge/conf_wb_err_pending_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_wb_err_pending_out )
    );
    X_OR2 \bridge/conf_wb_err_pending_out/FFY/ASYNC_FF_GSR_OR_154 (
      .I0 (\bridge/configuration/delete_wb_err_cs_bit8 ),
      .I1 (GSR),
      .O (\bridge/conf_wb_err_pending_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_ba0_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_ba0_out[13]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<24> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N34 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba0_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba0_out [12])
    );
    X_OR2 \bridge/conf_pci_ba0_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba0_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba0_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<25> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N34 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba0_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba0_out [13])
    );
    X_OR2 \bridge/conf_pci_ba0_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba0_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba0_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr0<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr0[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N79 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [16])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N79 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [17])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_base_addr0<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_base_addr0[19]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N79 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [18])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N79 ),
      .SET (GND),
      .RST (\bridge/configuration/pci_base_addr0[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_base_addr0 [19])
    );
    X_OR2 \bridge/configuration/pci_base_addr0<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_base_addr0[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_base_addr0[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_ba0_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_ba0_out[15]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<26> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N34 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba0_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba0_out [14])
    );
    X_OR2 \bridge/conf_pci_ba0_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba0_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba0_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<27> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N34 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba0_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba0_out [15])
    );
    X_OR2 \bridge/conf_pci_ba0_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba0_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba0_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<10> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [10]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [10])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<11> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [11]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [11])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[11]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/conf_pci_ba0_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_ba0_out[17]/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<28> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N34 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba0_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba0_out [16])
    );
    X_OR2 \bridge/conf_pci_ba0_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba0_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba0_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_ba0_bit31_12_reg<29> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C285/N34 ),
      .SET (GND),
      .RST (\bridge/conf_pci_ba0_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_ba0_out [17])
    );
    X_OR2 \bridge/conf_pci_ba0_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_pci_ba0_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_ba0_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<20> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [20])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<21> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [21])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[21]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<12> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [12])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<13> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [13])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[13]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<30> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [30])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<31> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [31])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[31]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<22> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [22])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<23> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [23])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[23]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<14> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [14])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<15> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [15])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[15]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbr_waddr<0>/BYMUX (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_waddr [0]),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/BYNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/waddr_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST (\bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr [0])
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbr_waddr<0>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/FFY/RST )
    );
    X_OR2 \bridge/wishbone_slave_unit/fifos/wbr_waddr<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_waddr[0]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<24> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [24])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<25> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [25])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[25]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<16> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [16])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<17> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [17])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[17]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<26> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [26])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<27> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [27])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[27]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<18> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [18])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<19> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [19])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[19]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<28> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [28])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg_reg<29> (
      .I (\bridge/pci_target_unit/fifos_pcir_data_out [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_load_medium_reg_out ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg [29])
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/pcir_fifo_data_reg[29]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/configuration/pci_err_addr<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[1]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<0> (
      .I (\bridge/pciu_err_addr_out[0] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [0])
    );
    X_OR2 \bridge/configuration/pci_err_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<1> (
      .I (\bridge/pciu_err_addr_out[1] ),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [1])
    );
    X_OR2 \bridge/configuration/pci_err_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[3]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<2> (
      .I (ADR_O[2]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [2])
    );
    X_OR2 \bridge/configuration/pci_err_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<3> (
      .I (ADR_O[3]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [3])
    );
    X_OR2 \bridge/configuration/pci_err_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[5]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<4> (
      .I (ADR_O[4]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [4])
    );
    X_OR2 \bridge/configuration/pci_err_addr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<5> (
      .I (ADR_O[5]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [5])
    );
    X_OR2 \bridge/configuration/pci_err_addr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_ONE \bridge/configuration/status_bit15_11<14>/LOGIC_ONE (
      .O (\bridge/configuration/status_bit15_11[14]/LOGIC_ONE )
    );
    X_FF \bridge/configuration/status_bit15_11_reg2<14> (
      .I (\bridge/configuration/status_bit15_11[14]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/parchk_sig_serr_out ),
      .SET (GND),
      .RST (\bridge/configuration/status_bit15_11[14]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/status_bit15_11 [14])
    );
    X_OR2 \bridge/configuration/status_bit15_11<14>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/delete_status_bit14 ),
      .I1 (GSR),
      .O (\bridge/configuration/status_bit15_11[14]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[7]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<6> (
      .I (ADR_O[6]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [6])
    );
    X_OR2 \bridge/configuration/pci_err_addr<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<7> (
      .I (ADR_O[7]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [7])
    );
    X_OR2 \bridge/configuration/pci_err_addr<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/configuration/pci_err_addr<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/configuration/pci_err_addr[9]/SRNOT )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<8> (
      .I (ADR_O[8]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [8])
    );
    X_OR2 \bridge/configuration/pci_err_addr<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/pci_err_addr_reg<9> (
      .I (ADR_O[9]),
      .CLK (CLK_BUFGPed),
      .CE (N12311),
      .SET (GND),
      .RST (\bridge/configuration/pci_err_addr[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_err_addr [9])
    );
    X_OR2 \bridge/configuration/pci_err_addr<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/pci_err_addr[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_err_addr[9]/FFX/ASYNC_FF_GSR_OR )
    );
    X_ONE \bridge/configuration/status_bit15_11<13>/LOGIC_ONE (
      .O (\bridge/configuration/status_bit15_11[13]/LOGIC_ONE )
    );
    X_FF \bridge/configuration/status_bit15_11_reg3<13> (
      .I (\bridge/configuration/status_bit15_11[13]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wbu_mabort_rec_out ),
      .SET (GND),
      .RST (\bridge/configuration/status_bit15_11[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/status_bit15_11 [13])
    );
    X_OR2 \bridge/configuration/status_bit15_11<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/delete_status_bit13 ),
      .I1 (GSR),
      .O (\bridge/configuration/status_bit15_11[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_ONE \bridge/configuration/status_bit15_11<12>/LOGIC_ONE (
      .O (\bridge/configuration/status_bit15_11[12]/LOGIC_ONE )
    );
    X_FF \bridge/configuration/status_bit15_11_reg4<12> (
      .I (\bridge/configuration/status_bit15_11[12]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_sm_mabort_out ),
      .SET (GND),
      .RST (\bridge/configuration/status_bit15_11[12]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/status_bit15_11 [12])
    );
    X_OR2 \bridge/configuration/status_bit15_11<12>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/delete_status_bit12 ),
      .I1 (GSR),
      .O (\bridge/configuration/status_bit15_11[12]/FFY/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[11]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<10> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [10]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [10])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<11> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [11]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [11])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[11]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [0])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<1>/FFY/SETOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFY/SET )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFY/SET ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [1])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<1>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[21]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<20> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [20]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [20])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<21> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [21]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [21])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[13]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<12> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [12]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [12])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<13> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [13]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [13])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [2])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<3>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [3])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<3>/FFX/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFX/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[31]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<30> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [30]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [30])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<31> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [31]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [31])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[23]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<22> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [22]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [22])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<23> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [23]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [23])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[15]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<14> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [14]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [14])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<15> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [15]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [15])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [4])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<5>/FFY/RSTOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFY/RST )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr_reg<5> (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_next [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFX/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr [5])
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<5>/FFX/SETOR (
      .I (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/clear ),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFX/SET )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFX/SET ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbr_fifo_ctrl/wgrey_addr[5]/FFX/ASYNC_FF_GSR_OR )

    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[25]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<24> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [24]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [24])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<25> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [25]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [25])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[17]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<16> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [16]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [16])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<17> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [17]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [17])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/conf_pci_mem_io1_out/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_pci_mem_io1_out/SRNOT )
    );
    X_FF \bridge/configuration/pci_ba1_bit0_reg (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C287/N3 ),
      .SET (GND),
      .RST (\bridge/conf_pci_mem_io1_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_pci_mem_io1_out )
    );
    X_OR2 \bridge/conf_pci_mem_io1_out/FFY/ASYNC_FF_GSR_OR_155 (
      .I0 (\bridge/conf_pci_mem_io1_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_pci_mem_io1_out/FFY/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/C1140 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1140 (
      .ADR0 (\bridge/out_bckp_cbe_out [2]),
      .ADR1 (\bridge/out_bckp_cbe_out [1]),
      .ADR2 (\bridge/out_bckp_cbe_out [0]),
      .ADR3 (\bridge/out_bckp_cbe_out [3]),
      .O (\bridge/parity_checker/BLK0_4/GROM )
    );
    defparam \bridge/parity_checker/C1125 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1125 (
      .ADR0 (\bridge/parity_checker/syn3204 ),
      .ADR1 (\bridge/parity_checker/syn3210 ),
      .ADR2 (\bridge/parity_checker/par_cbe_out ),
      .ADR3 (\bridge/parity_checker/syn3125 ),
      .O (\bridge/parity_checker/syn3234 )
    );
    X_XOR2 \bridge/parity_checker/C1124 (
      .I0 (\bridge/parity_checker/syn3214 ),
      .I1 (\bridge/parity_checker/syn3234 ),
      .O (\bridge/parity_checker/BLK0_4/XORF )
    );
    X_BUF \bridge/parity_checker/BLK0_4/YUSED (
      .I (\bridge/parity_checker/BLK0_4/GROM ),
      .O (\bridge/parity_checker/par_cbe_out )
    );
    X_BUF \bridge/parity_checker/BLK0_4/XUSED (
      .I (\bridge/parity_checker/BLK0_4/XORF ),
      .O (\bridge/parity_checker/par_out_only )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<11>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[11]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<10> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [10]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [10])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<11> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [11]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [11])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[11]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/C1129 .INIT = 16'h9966;
    X_LUT4 \bridge/parity_checker/C1129 (
      .ADR0 (\bridge/out_bckp_ad_out [16]),
      .ADR1 (\bridge/out_bckp_ad_out [3]),
      .ADR2 (VCC),
      .ADR3 (\bridge/out_bckp_ad_out [2]),
      .O (\bridge/parity_checker/BLK1_4/GROM )
    );
    defparam \bridge/parity_checker/C1128 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1128 (
      .ADR0 (\bridge/out_bckp_ad_out [10]),
      .ADR1 (\bridge/parity_checker/syn3190 ),
      .ADR2 (\bridge/parity_checker/syn3208 ),
      .ADR3 (\bridge/parity_checker/syn3189 ),
      .O (\bridge/parity_checker/syn3232 )
    );
    X_XOR2 \bridge/parity_checker/C1127 (
      .I0 (\bridge/parity_checker/BLK1_4/CYINIT ),
      .I1 (\bridge/parity_checker/syn3232 ),
      .O (\bridge/parity_checker/BLK1_4/XORF )
    );
    X_BUF \bridge/parity_checker/BLK1_4/CYINIT_156 (
      .I (\bridge/out_bckp_ad_out [15]),
      .O (\bridge/parity_checker/BLK1_4/CYINIT )
    );
    X_BUF \bridge/parity_checker/BLK1_4/YUSED (
      .I (\bridge/parity_checker/BLK1_4/GROM ),
      .O (\bridge/parity_checker/syn3208 )
    );
    X_BUF \bridge/parity_checker/BLK1_4/XUSED (
      .I (\bridge/parity_checker/BLK1_4/XORF ),
      .O (\bridge/parity_checker/syn3210 )
    );
    defparam \bridge/parity_checker/C1134 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1134 (
      .ADR0 (\bridge/out_bckp_ad_out [24]),
      .ADR1 (\bridge/out_bckp_ad_out [26]),
      .ADR2 (\bridge/out_bckp_ad_out [25]),
      .ADR3 (\bridge/out_bckp_ad_out [27]),
      .O (\bridge/parity_checker/BLK2_4/GROM )
    );
    defparam \bridge/parity_checker/C1133 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1133 (
      .ADR0 (\bridge/out_bckp_ad_out [28]),
      .ADR1 (\bridge/out_bckp_ad_out [29]),
      .ADR2 (\bridge/parity_checker/syn3196 ),
      .ADR3 (\bridge/out_bckp_ad_out [30]),
      .O (\bridge/parity_checker/syn3230 )
    );
    X_XOR2 \bridge/parity_checker/C1132 (
      .I0 (\bridge/parity_checker/BLK2_4/CYINIT ),
      .I1 (\bridge/parity_checker/syn3230 ),
      .O (\bridge/parity_checker/BLK2_4/XORF )
    );
    X_BUF \bridge/parity_checker/BLK2_4/CYINIT_157 (
      .I (\bridge/out_bckp_ad_out [31]),
      .O (\bridge/parity_checker/BLK2_4/CYINIT )
    );
    X_BUF \bridge/parity_checker/BLK2_4/YUSED (
      .I (\bridge/parity_checker/BLK2_4/GROM ),
      .O (\bridge/parity_checker/syn3196 )
    );
    X_BUF \bridge/parity_checker/BLK2_4/XUSED (
      .I (\bridge/parity_checker/BLK2_4/XORF ),
      .O (\bridge/parity_checker/syn3125 )
    );
    X_ONE \bridge/configuration/status_bit15_11<11>/LOGIC_ONE (
      .O (\bridge/configuration/status_bit15_11[11]/LOGIC_ONE )
    );
    X_FF \bridge/configuration/status_bit15_11_reg5<11> (
      .I (\bridge/configuration/status_bit15_11[11]/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pciu_pciif_tabort_set_out ),
      .SET (GND),
      .RST (\bridge/configuration/status_bit15_11[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/status_bit15_11 [11])
    );
    X_OR2 \bridge/configuration/status_bit15_11<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/configuration/delete_status_bit11 ),
      .I1 (GSR),
      .O (\bridge/configuration/status_bit15_11[11]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C17944.INIT = 16'h9009;
    X_LUT4 C17944(
      .ADR0 (\bridge/pci_target_unit/del_sync_addr_out [6]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .ADR3 (\bridge/pci_target_unit/del_sync_addr_out [7]),
      .O (\bridge/parity_checker/BLK3_4/GROM )
    );
    defparam \bridge/parity_checker/C1144 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1144 (
      .ADR0 (\bridge/parity_checker/cbe_par_reg ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .O (\bridge/parity_checker/syn3228 )
    );
    X_XOR2 \bridge/parity_checker/C1143 (
      .I0 (\bridge/parity_checker/syn3172 ),
      .I1 (\bridge/parity_checker/syn3228 ),
      .O (\bridge/parity_checker/BLK3_4/XORF )
    );
    X_BUF \bridge/parity_checker/BLK3_4/YUSED (
      .I (\bridge/parity_checker/BLK3_4/GROM ),
      .O (syn182000)
    );
    X_BUF \bridge/parity_checker/BLK3_4/XUSED (
      .I (\bridge/parity_checker/BLK3_4/XORF ),
      .O (\bridge/parity_checker/syn3174 )
    );
    defparam \bridge/parity_checker/C1148 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1148 (
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .O (\bridge/parity_checker/BLK4_4/GROM )
    );
    defparam \bridge/parity_checker/C1147 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/C1147 (
      .ADR0 (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .ADR2 (\bridge/parity_checker/syn3148 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .O (\bridge/parity_checker/syn3226 )
    );
    X_XOR2 \bridge/parity_checker/C1146 (
      .I0 (\bridge/parity_checker/BLK4_4/CYINIT ),
      .I1 (\bridge/parity_checker/syn3226 ),
      .O (\bridge/parity_checker/BLK4_4/XORF )
    );
    X_BUF \bridge/parity_checker/BLK4_4/CYINIT_158 (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .O (\bridge/parity_checker/BLK4_4/CYINIT )
    );
    X_BUF \bridge/parity_checker/BLK4_4/YUSED (
      .I (\bridge/parity_checker/BLK4_4/GROM ),
      .O (\bridge/parity_checker/syn3148 )
    );
    X_BUF \bridge/parity_checker/BLK4_4/XUSED (
      .I (\bridge/parity_checker/BLK4_4/XORF ),
      .O (\bridge/parity_checker/syn3083 )
    );
    X_INV \CRT/pix_start_addr<11>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[11]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<10> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [10]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[11]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [10])
    );
    X_OR2 \CRT/pix_start_addr<11>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[11]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[11]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<11> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [11]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[11]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [11])
    );
    X_OR2 \CRT/pix_start_addr<11>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[11]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[11]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/parity_checker/par_gen/C74 .INIT = 16'h6996;
    X_LUT4 \bridge/parity_checker/par_gen/C74 (
      .ADR0 (N_CBE[3]),
      .ADR1 (N_CBE[2]),
      .ADR2 (N_CBE[0]),
      .ADR3 (N_CBE[1]),
      .O (\bridge/parity_checker/par_gen/syn156 )
    );
    X_XOR2 \bridge/parity_checker/par_gen/C73 (
      .I0 (\bridge/parity_checker/data_par ),
      .I1 (\bridge/parity_checker/par_gen/syn156 ),
      .O (\bridge/parity_checker/par_gen/BLK0_2/XORF )
    );
    X_BUF \bridge/parity_checker/par_gen/BLK0_2/XUSED (
      .I (\bridge/parity_checker/par_gen/BLK0_2/XORF ),
      .O (\bridge/parity_checker/par_gen/syn143 )
    );
    X_BUF \C15440/IBUF (
      .I (RST),
      .O (\RST/IBUF )
    );
    X_KEEPER \RST/KEEPER_159 (
      .O (\RST/KEEPER )
    );
    X_IPAD \RST/PAD (
      .PAD (RST)
    );
    X_BUF \RST/IMUX (
      .I (\RST/IBUF ),
      .O (N_RST)
    );
    X_BUF \AD<27>/DELAY (
      .I (N_AD[27]),
      .O (\AD[27]/IDELAY )
    );
    X_BUF \C15406/IBUF (
      .I (AD[27]),
      .O (N_AD[27])
    );
    X_INV \AD<27>/ENABLEINV (
      .I (AD_en[27]),
      .O (\AD[27]/ENABLE )
    );
    X_TRI \C15406/OBUFT (
      .I (AD_out[27]),
      .O (AD[27]),
      .CTL (\AD[27]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<27>/KEEPER (
      .O (\AD[27]/KEEPER )
    );
    X_BPAD \AD<27>/PAD (
      .PAD (AD[27])
    );
    X_INV \AD<27>/SRMUX (
      .I (N_RST),
      .O (\AD[27]/SRNOT )
    );
    X_BUF \AD<27>/OMUX (
      .I (\bridge/output_backup/C3/N168 ),
      .O (\AD[27]/OD )
    );
    X_AND2 \AD<27>/OUTBUF_GTS_AND (
      .I0 (\AD[27]/ENABLE ),
      .I1 (\AD[27]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[27]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<27> (
      .I (\AD[27]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[27]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [27])
    );
    X_OR2 \AD<27>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[27]/SRNOT ),
      .I1 (GSR),
      .O (\AD[27]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob27/dat_out_reg (
      .I (\AD[27]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_high ),
      .SET (GND),
      .RST (\AD[27]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[27])
    );
    X_OR2 \AD<27>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[27]/SRNOT ),
      .I1 (GSR),
      .O (\AD[27]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob27/en_out_reg (
      .I (N12338),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[27]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[27])
    );
    X_OR2 \AD<27>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[27]/SRNOT ),
      .I1 (GSR),
      .O (\AD[27]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<26>/DELAY (
      .I (N_AD[26]),
      .O (\AD[26]/IDELAY )
    );
    X_BUF \C15407/IBUF (
      .I (AD[26]),
      .O (N_AD[26])
    );
    X_INV \AD<26>/ENABLEINV (
      .I (AD_en[26]),
      .O (\AD[26]/ENABLE )
    );
    X_TRI \C15407/OBUFT (
      .I (AD_out[26]),
      .O (AD[26]),
      .CTL (\AD[26]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<26>/KEEPER (
      .O (\AD[26]/KEEPER )
    );
    X_BPAD \AD<26>/PAD (
      .PAD (AD[26])
    );
    X_INV \AD<26>/SRMUX (
      .I (N_RST),
      .O (\AD[26]/SRNOT )
    );
    X_BUF \AD<26>/OMUX (
      .I (\bridge/output_backup/C3/N162 ),
      .O (\AD[26]/OD )
    );
    X_AND2 \AD<26>/OUTBUF_GTS_AND (
      .I0 (\AD[26]/ENABLE ),
      .I1 (\AD[26]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[26]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<26> (
      .I (\AD[26]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[26]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [26])
    );
    X_OR2 \AD<26>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[26]/SRNOT ),
      .I1 (GSR),
      .O (\AD[26]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob26/dat_out_reg (
      .I (\AD[26]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_high ),
      .SET (GND),
      .RST (\AD[26]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[26])
    );
    X_OR2 \AD<26>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[26]/SRNOT ),
      .I1 (GSR),
      .O (\AD[26]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob26/en_out_reg (
      .I (N12338),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[26]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[26])
    );
    X_OR2 \AD<26>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[26]/SRNOT ),
      .I1 (GSR),
      .O (\AD[26]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<25>/DELAY (
      .I (N_AD[25]),
      .O (\AD[25]/IDELAY )
    );
    X_BUF \C15408/IBUF (
      .I (AD[25]),
      .O (N_AD[25])
    );
    X_INV \AD<25>/ENABLEINV (
      .I (AD_en[25]),
      .O (\AD[25]/ENABLE )
    );
    X_TRI \C15408/OBUFT (
      .I (AD_out[25]),
      .O (AD[25]),
      .CTL (\AD[25]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<25>/KEEPER (
      .O (\AD[25]/KEEPER )
    );
    X_BPAD \AD<25>/PAD (
      .PAD (AD[25])
    );
    X_INV \AD<25>/SRMUX (
      .I (N_RST),
      .O (\AD[25]/SRNOT )
    );
    X_BUF \AD<25>/OMUX (
      .I (\bridge/output_backup/C3/N156 ),
      .O (\AD[25]/OD )
    );
    X_AND2 \AD<25>/OUTBUF_GTS_AND (
      .I0 (\AD[25]/ENABLE ),
      .I1 (\AD[25]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[25]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<25> (
      .I (\AD[25]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[25]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [25])
    );
    X_OR2 \AD<25>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[25]/SRNOT ),
      .I1 (GSR),
      .O (\AD[25]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob25/dat_out_reg (
      .I (\AD[25]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_high ),
      .SET (GND),
      .RST (\AD[25]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[25])
    );
    X_OR2 \AD<25>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[25]/SRNOT ),
      .I1 (GSR),
      .O (\AD[25]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob25/en_out_reg (
      .I (N12338),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[25]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[25])
    );
    X_OR2 \AD<25>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[25]/SRNOT ),
      .I1 (GSR),
      .O (\AD[25]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<24>/DELAY (
      .I (N_AD[24]),
      .O (\AD[24]/IDELAY )
    );
    X_BUF \C15409/IBUF (
      .I (AD[24]),
      .O (N_AD[24])
    );
    X_INV \AD<24>/ENABLEINV (
      .I (AD_en[24]),
      .O (\AD[24]/ENABLE )
    );
    X_TRI \C15409/OBUFT (
      .I (AD_out[24]),
      .O (AD[24]),
      .CTL (\AD[24]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<24>/KEEPER (
      .O (\AD[24]/KEEPER )
    );
    X_BPAD \AD<24>/PAD (
      .PAD (AD[24])
    );
    X_INV \AD<24>/SRMUX (
      .I (N_RST),
      .O (\AD[24]/SRNOT )
    );
    X_BUF \AD<24>/OMUX (
      .I (\bridge/output_backup/C3/N150 ),
      .O (\AD[24]/OD )
    );
    X_AND2 \AD<24>/OUTBUF_GTS_AND (
      .I0 (\AD[24]/ENABLE ),
      .I1 (\AD[24]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[24]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<24> (
      .I (\AD[24]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[24]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [24])
    );
    X_OR2 \AD<24>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[24]/SRNOT ),
      .I1 (GSR),
      .O (\AD[24]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob24/dat_out_reg (
      .I (\AD[24]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_high ),
      .SET (GND),
      .RST (\AD[24]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[24])
    );
    X_OR2 \AD<24>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[24]/SRNOT ),
      .I1 (GSR),
      .O (\AD[24]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob24/en_out_reg (
      .I (N12338),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[24]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[24])
    );
    X_OR2 \AD<24>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[24]/SRNOT ),
      .I1 (GSR),
      .O (\AD[24]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<23>/DELAY (
      .I (N_AD[23]),
      .O (\AD[23]/IDELAY )
    );
    X_BUF \C15410/IBUF (
      .I (AD[23]),
      .O (N_AD[23])
    );
    X_INV \AD<23>/ENABLEINV (
      .I (AD_en[23]),
      .O (\AD[23]/ENABLE )
    );
    X_TRI \C15410/OBUFT (
      .I (AD_out[23]),
      .O (AD[23]),
      .CTL (\AD[23]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<23>/KEEPER (
      .O (\AD[23]/KEEPER )
    );
    X_BPAD \AD<23>/PAD (
      .PAD (AD[23])
    );
    X_INV \AD<23>/SRMUX (
      .I (N_RST),
      .O (\AD[23]/SRNOT )
    );
    X_BUF \AD<23>/OMUX (
      .I (\bridge/output_backup/C3/N144 ),
      .O (\AD[23]/OD )
    );
    X_AND2 \AD<23>/OUTBUF_GTS_AND (
      .I0 (\AD[23]/ENABLE ),
      .I1 (\AD[23]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[23]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<23> (
      .I (\AD[23]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[23]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [23])
    );
    X_OR2 \AD<23>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[23]/SRNOT ),
      .I1 (GSR),
      .O (\AD[23]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob23/dat_out_reg (
      .I (\AD[23]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mhigh ),
      .SET (GND),
      .RST (\AD[23]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[23])
    );
    X_OR2 \AD<23>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[23]/SRNOT ),
      .I1 (GSR),
      .O (\AD[23]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob23/en_out_reg (
      .I (N12330),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[23]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[23])
    );
    X_OR2 \AD<23>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[23]/SRNOT ),
      .I1 (GSR),
      .O (\AD[23]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \CBE<3>/DELAY (
      .I (\CBE[3]/IBUF ),
      .O (\CBE[3]/IDELAY )
    );
    X_BUF \C15434/IBUF (
      .I (CBE[3]),
      .O (\CBE[3]/IBUF )
    );
    X_INV \CBE<3>/ENABLEINV (
      .I (CBE_en[3]),
      .O (\CBE[3]/ENABLE )
    );
    X_TRI \C15434/OBUFT (
      .I (CBE_out[3]),
      .O (CBE[3]),
      .CTL (\CBE[3]/OUTBUF_GTS_AND )
    );
    X_KEEPER \CBE<3>/KEEPER (
      .O (\CBE[3]/KEEPER )
    );
    X_BPAD \CBE<3>/PAD (
      .PAD (CBE[3])
    );
    X_INV \CBE<3>/SRMUX (
      .I (N_RST),
      .O (\CBE[3]/SRNOT )
    );
    X_BUF \CBE<3>/IMUX (
      .I (\CBE[3]/IBUF ),
      .O (N_CBE[3])
    );
    X_BUF \CBE<3>/OMUX (
      .I (\bridge/pci_mux_cbe_in [3]),
      .O (\CBE[3]/OD )
    );
    X_INV \CBE<3>/TRIMUX (
      .I (\bridge/pci_mux_cbe_en_in ),
      .O (\CBE[3]/TNOT )
    );
    X_AND2 \CBE<3>/OUTBUF_GTS_AND (
      .I0 (\CBE[3]/ENABLE ),
      .I1 (\CBE[3]/OUTBUF_GTS_AND_1_INV ),
      .O (\CBE[3]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_cbe_reg_out_reg<3> (
      .I (\CBE[3]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CBE[3]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/in_reg_cbe_out [3])
    );
    X_OR2 \CBE<3>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[3]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[3]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/cbe_iob3/dat_out_reg (
      .I (\CBE[3]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_mas_load_in ),
      .SET (GND),
      .RST (\CBE[3]/OFF/ASYNC_FF_GSR_OR ),
      .O (CBE_out[3])
    );
    X_OR2 \CBE<3>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[3]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[3]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/cbe_iob3/en_out_reg (
      .I (\CBE[3]/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\CBE[3]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (CBE_en[3])
    );
    X_OR2 \CBE<3>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[3]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[3]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF C_IDSEL(
      .I (IDSEL),
      .O (\IDSEL/IBUF )
    );
    X_KEEPER \IDSEL/KEEPER_160 (
      .O (\IDSEL/KEEPER )
    );
    X_IPAD \IDSEL/PAD (
      .PAD (IDSEL)
    );
    X_BUF \IDSEL/IMUX (
      .I (\IDSEL/IBUF ),
      .O (N_IDSEL)
    );
    X_BUF \AD<17>/DELAY (
      .I (N_AD[17]),
      .O (\AD[17]/IDELAY )
    );
    X_BUF \C15416/IBUF (
      .I (AD[17]),
      .O (N_AD[17])
    );
    X_INV \AD<17>/ENABLEINV (
      .I (AD_en[17]),
      .O (\AD[17]/ENABLE )
    );
    X_TRI \C15416/OBUFT (
      .I (AD_out[17]),
      .O (AD[17]),
      .CTL (\AD[17]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<17>/KEEPER (
      .O (\AD[17]/KEEPER )
    );
    X_BPAD \AD<17>/PAD (
      .PAD (AD[17])
    );
    X_INV \AD<17>/SRMUX (
      .I (N_RST),
      .O (\AD[17]/SRNOT )
    );
    X_AND2 \AD<17>/OUTBUF_GTS_AND (
      .I0 (\AD[17]/ENABLE ),
      .I1 (\AD[17]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[17]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<17> (
      .I (\AD[17]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[17]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [17])
    );
    X_OR2 \AD<17>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[17]/SRNOT ),
      .I1 (GSR),
      .O (\AD[17]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob17/dat_out_reg (
      .I (\bridge/output_backup/C3/N108 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mhigh ),
      .SET (GND),
      .RST (\AD[17]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[17])
    );
    X_OR2 \AD<17>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[17]/SRNOT ),
      .I1 (GSR),
      .O (\AD[17]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob17/en_out_reg (
      .I (N12330),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[17]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[17])
    );
    X_OR2 \AD<17>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[17]/SRNOT ),
      .I1 (GSR),
      .O (\AD[17]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<16>/DELAY (
      .I (N_AD[16]),
      .O (\AD[16]/IDELAY )
    );
    X_BUF \C15417/IBUF (
      .I (AD[16]),
      .O (N_AD[16])
    );
    X_INV \AD<16>/ENABLEINV (
      .I (AD_en[16]),
      .O (\AD[16]/ENABLE )
    );
    X_TRI \C15417/OBUFT (
      .I (AD_out[16]),
      .O (AD[16]),
      .CTL (\AD[16]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<16>/KEEPER (
      .O (\AD[16]/KEEPER )
    );
    X_BPAD \AD<16>/PAD (
      .PAD (AD[16])
    );
    X_INV \AD<16>/SRMUX (
      .I (N_RST),
      .O (\AD[16]/SRNOT )
    );
    X_BUF \AD<16>/OMUX (
      .I (\bridge/output_backup/C3/N102 ),
      .O (\AD[16]/OD )
    );
    X_AND2 \AD<16>/OUTBUF_GTS_AND (
      .I0 (\AD[16]/ENABLE ),
      .I1 (\AD[16]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[16]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<16> (
      .I (\AD[16]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[16]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [16])
    );
    X_OR2 \AD<16>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[16]/SRNOT ),
      .I1 (GSR),
      .O (\AD[16]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob16/dat_out_reg (
      .I (\AD[16]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mhigh ),
      .SET (GND),
      .RST (\AD[16]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[16])
    );
    X_OR2 \AD<16>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[16]/SRNOT ),
      .I1 (GSR),
      .O (\AD[16]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob16/en_out_reg (
      .I (N12330),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[16]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[16])
    );
    X_OR2 \AD<16>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[16]/SRNOT ),
      .I1 (GSR),
      .O (\AD[16]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \CBE<2>/DELAY (
      .I (\CBE[2]/IBUF ),
      .O (\CBE[2]/IDELAY )
    );
    X_BUF \C15435/IBUF (
      .I (CBE[2]),
      .O (\CBE[2]/IBUF )
    );
    X_INV \CBE<2>/ENABLEINV (
      .I (CBE_en[2]),
      .O (\CBE[2]/ENABLE )
    );
    X_TRI \C15435/OBUFT (
      .I (CBE_out[2]),
      .O (CBE[2]),
      .CTL (\CBE[2]/OUTBUF_GTS_AND )
    );
    X_KEEPER \CBE<2>/KEEPER (
      .O (\CBE[2]/KEEPER )
    );
    X_BPAD \CBE<2>/PAD (
      .PAD (CBE[2])
    );
    X_INV \CBE<2>/SRMUX (
      .I (N_RST),
      .O (\CBE[2]/SRNOT )
    );
    X_BUF \CBE<2>/IMUX (
      .I (\CBE[2]/IBUF ),
      .O (N_CBE[2])
    );
    X_BUF \CBE<2>/OMUX (
      .I (\bridge/pci_mux_cbe_in [2]),
      .O (\CBE[2]/OD )
    );
    X_INV \CBE<2>/TRIMUX (
      .I (\bridge/pci_mux_cbe_en_in ),
      .O (\CBE[2]/TNOT )
    );
    X_AND2 \CBE<2>/OUTBUF_GTS_AND (
      .I0 (\CBE[2]/ENABLE ),
      .I1 (\CBE[2]/OUTBUF_GTS_AND_1_INV ),
      .O (\CBE[2]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_cbe_reg_out_reg<2> (
      .I (\CBE[2]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CBE[2]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/in_reg_cbe_out [2])
    );
    X_OR2 \CBE<2>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[2]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[2]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/cbe_iob2/dat_out_reg (
      .I (\CBE[2]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_mas_load_in ),
      .SET (GND),
      .RST (\CBE[2]/OFF/ASYNC_FF_GSR_OR ),
      .O (CBE_out[2])
    );
    X_OR2 \CBE<2>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[2]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[2]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/cbe_iob2/en_out_reg (
      .I (\CBE[2]/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\CBE[2]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (CBE_en[2])
    );
    X_OR2 \CBE<2>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[2]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[2]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[27]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<26> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [26]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [26])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<27> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [27]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [27])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \STOP/DELAY (
      .I (\STOP/IBUF ),
      .O (\STOP/IDELAY )
    );
    X_BUF \C15450/IBUF (
      .I (STOP),
      .O (\STOP/IBUF )
    );
    X_INV \STOP/ENABLEINV (
      .I (STOP_en),
      .O (\STOP/ENABLE )
    );
    X_TRI \C15450/OBUFT (
      .I (STOP_out),
      .O (STOP),
      .CTL (\STOP/OUTBUF_GTS_AND )
    );
    X_KEEPER \STOP/KEEPER_161 (
      .O (\STOP/KEEPER )
    );
    X_BPAD \STOP/PAD (
      .PAD (STOP)
    );
    X_INV \STOP/SRMUX (
      .I (N_RST),
      .O (\STOP/SRNOT )
    );
    X_BUF \STOP/IMUX (
      .I (\STOP/IBUF ),
      .O (N_STOP)
    );
    X_INV \STOP/TRIMUX (
      .I (\bridge/pciu_pciif_devsel_en_out ),
      .O (\STOP/TNOT )
    );
    X_AND2 \STOP/OUTBUF_GTS_AND_162 (
      .I0 (\STOP/ENABLE ),
      .I1 (\STOP/OUTBUF_GTS_AND_1_INV ),
      .O (\STOP/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_stop_reg_out_reg (
      .I (\STOP/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\STOP/IFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/in_reg_stop_out )
    );
    X_OR2 \STOP/IFF/ASYNC_FF_GSR_OR_163 (
      .I0 (\STOP/SRNOT ),
      .I1 (GSR),
      .O (\STOP/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/stop_iob/dat_out_reg (
      .I (N12476),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\STOP/OFF/ASYNC_FF_GSR_OR ),
      .O (STOP_out)
    );
    X_OR2 \STOP/OFF/ASYNC_FF_GSR_OR_164 (
      .I0 (\STOP/SRNOT ),
      .I1 (GSR),
      .O (\STOP/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/stop_iob/en_out_reg (
      .I (\STOP/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\STOP/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (STOP_en)
    );
    X_OR2 \STOP/TFF/ASYNC_FF_GSR_OR_165 (
      .I0 (\STOP/SRNOT ),
      .I1 (GSR),
      .O (\STOP/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<22>/DELAY (
      .I (N_AD[22]),
      .O (\AD[22]/IDELAY )
    );
    X_BUF \C15411/IBUF (
      .I (AD[22]),
      .O (N_AD[22])
    );
    X_INV \AD<22>/ENABLEINV (
      .I (AD_en[22]),
      .O (\AD[22]/ENABLE )
    );
    X_TRI \C15411/OBUFT (
      .I (AD_out[22]),
      .O (AD[22]),
      .CTL (\AD[22]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<22>/KEEPER (
      .O (\AD[22]/KEEPER )
    );
    X_BPAD \AD<22>/PAD (
      .PAD (AD[22])
    );
    X_INV \AD<22>/SRMUX (
      .I (N_RST),
      .O (\AD[22]/SRNOT )
    );
    X_BUF \AD<22>/OMUX (
      .I (\bridge/output_backup/C3/N138 ),
      .O (\AD[22]/OD )
    );
    X_AND2 \AD<22>/OUTBUF_GTS_AND (
      .I0 (\AD[22]/ENABLE ),
      .I1 (\AD[22]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[22]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<22> (
      .I (\AD[22]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[22]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [22])
    );
    X_OR2 \AD<22>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[22]/SRNOT ),
      .I1 (GSR),
      .O (\AD[22]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob22/dat_out_reg (
      .I (\AD[22]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mhigh ),
      .SET (GND),
      .RST (\AD[22]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[22])
    );
    X_OR2 \AD<22>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[22]/SRNOT ),
      .I1 (GSR),
      .O (\AD[22]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob22/en_out_reg (
      .I (N12330),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[22]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[22])
    );
    X_OR2 \AD<22>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[22]/SRNOT ),
      .I1 (GSR),
      .O (\AD[22]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[19]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<18> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [18]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [18])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<19> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [19]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [19])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \FRAME/DELAY (
      .I (\FRAME/IBUF ),
      .O (\FRAME/IDELAY )
    );
    X_BUF \C15445/IBUF (
      .I (FRAME),
      .O (\FRAME/IBUF )
    );
    X_INV \FRAME/ENABLEINV (
      .I (FRAME_en),
      .O (\FRAME/ENABLE )
    );
    X_TRI \C15445/OBUFT (
      .I (FRAME_out),
      .O (FRAME),
      .CTL (\FRAME/OUTBUF_GTS_AND )
    );
    X_KEEPER \FRAME/KEEPER_166 (
      .O (\FRAME/KEEPER )
    );
    X_BPAD \FRAME/PAD (
      .PAD (FRAME)
    );
    X_INV \FRAME/SRMUX (
      .I (N_RST),
      .O (\FRAME/SRNOT )
    );
    X_BUF \FRAME/IMUX (
      .I (\FRAME/IBUF ),
      .O (N_FRAME)
    );
    X_INV \FRAME/TRIMUX (
      .I (\bridge/pci_mux_frame_en_in ),
      .O (\FRAME/TNOT )
    );
    X_AND2 \FRAME/OUTBUF_GTS_AND_167 (
      .I0 (\FRAME/ENABLE ),
      .I1 (\FRAME/OUTBUF_GTS_AND_1_INV ),
      .O (\FRAME/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_frame_reg_out_reg (
      .I (\FRAME/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\FRAME/IFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/in_reg_frame_out )
    );
    X_OR2 \FRAME/IFF/ASYNC_FF_GSR_OR_168 (
      .I0 (\FRAME/SRNOT ),
      .I1 (GSR),
      .O (\FRAME/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/frame_iob/dat_out_reg (
      .I (\bridge/pci_mux_frame_in ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_frame_load_in ),
      .SET (GND),
      .RST (\FRAME/OFF/ASYNC_FF_GSR_OR ),
      .O (FRAME_out)
    );
    X_OR2 \FRAME/OFF/ASYNC_FF_GSR_OR_169 (
      .I0 (\FRAME/SRNOT ),
      .I1 (GSR),
      .O (\FRAME/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/frame_iob/en_out_reg (
      .I (\FRAME/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\FRAME/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (FRAME_en)
    );
    X_OR2 \FRAME/TFF/ASYNC_FF_GSR_OR_170 (
      .I0 (\FRAME/SRNOT ),
      .I1 (GSR),
      .O (\FRAME/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \C15452/IBUF (
      .I (PERR),
      .O (\PERR/IBUF )
    );
    X_INV \PERR/ENABLEINV (
      .I (PERR_en),
      .O (\PERR/ENABLE )
    );
    X_TRI \C15452/OBUFT (
      .I (PERR_out),
      .O (PERR),
      .CTL (\PERR/OUTBUF_GTS_AND )
    );
    X_KEEPER \PERR/KEEPER_171 (
      .O (\PERR/KEEPER )
    );
    X_BPAD \PERR/PAD (
      .PAD (PERR)
    );
    X_INV \PERR/SRMUX (
      .I (N_RST),
      .O (\PERR/SRNOT )
    );
    X_BUF \PERR/IMUX (
      .I (\PERR/IBUF ),
      .O (N_PERR)
    );
    X_BUF \PERR/OMUX (
      .I (N12031),
      .O (\PERR/OD )
    );
    X_AND2 \PERR/OUTBUF_GTS_AND_172 (
      .I0 (\PERR/ENABLE ),
      .I1 (\PERR/OUTBUF_GTS_AND_1_INV ),
      .O (\PERR/OUTBUF_GTS_AND )
    );
    X_FF \bridge/pci_io_mux/perr_iob/dat_out_reg (
      .I (\PERR/OD ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\PERR/OFF/ASYNC_FF_GSR_OR ),
      .O (PERR_out)
    );
    X_OR2 \PERR/OFF/ASYNC_FF_GSR_OR_173 (
      .I0 (\PERR/SRNOT ),
      .I1 (GSR),
      .O (\PERR/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/perr_iob/en_out_reg (
      .I (N12033),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\PERR/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (PERR_en)
    );
    X_OR2 \PERR/TFF/ASYNC_FF_GSR_OR_174 (
      .I0 (\PERR/SRNOT ),
      .I1 (GSR),
      .O (\PERR/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<21>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[21]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<20> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [20]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [20])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<21> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [21]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [21])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[21]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<21>/DELAY (
      .I (N_AD[21]),
      .O (\AD[21]/IDELAY )
    );
    X_BUF \C15412/IBUF (
      .I (AD[21]),
      .O (N_AD[21])
    );
    X_INV \AD<21>/ENABLEINV (
      .I (AD_en[21]),
      .O (\AD[21]/ENABLE )
    );
    X_TRI \C15412/OBUFT (
      .I (AD_out[21]),
      .O (AD[21]),
      .CTL (\AD[21]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<21>/KEEPER (
      .O (\AD[21]/KEEPER )
    );
    X_BPAD \AD<21>/PAD (
      .PAD (AD[21])
    );
    X_INV \AD<21>/SRMUX (
      .I (N_RST),
      .O (\AD[21]/SRNOT )
    );
    X_BUF \AD<21>/OMUX (
      .I (\bridge/output_backup/C3/N132 ),
      .O (\AD[21]/OD )
    );
    X_AND2 \AD<21>/OUTBUF_GTS_AND (
      .I0 (\AD[21]/ENABLE ),
      .I1 (\AD[21]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[21]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<21> (
      .I (\AD[21]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[21]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [21])
    );
    X_OR2 \AD<21>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[21]/SRNOT ),
      .I1 (GSR),
      .O (\AD[21]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob21/dat_out_reg (
      .I (\AD[21]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mhigh ),
      .SET (GND),
      .RST (\AD[21]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[21])
    );
    X_OR2 \AD<21>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[21]/SRNOT ),
      .I1 (GSR),
      .O (\AD[21]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob21/en_out_reg (
      .I (N12330),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[21]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[21])
    );
    X_OR2 \AD<21>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[21]/SRNOT ),
      .I1 (GSR),
      .O (\AD[21]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \IRDY/DELAY (
      .I (\IRDY/IBUF ),
      .O (\IRDY/IDELAY )
    );
    X_BUF \C15446/IBUF (
      .I (IRDY),
      .O (\IRDY/IBUF )
    );
    X_INV \IRDY/ENABLEINV (
      .I (IRDY_en),
      .O (\IRDY/ENABLE )
    );
    X_TRI \C15446/OBUFT (
      .I (IRDY_out),
      .O (IRDY),
      .CTL (\IRDY/OUTBUF_GTS_AND )
    );
    X_KEEPER \IRDY/KEEPER_175 (
      .O (\IRDY/KEEPER )
    );
    X_BPAD \IRDY/PAD (
      .PAD (IRDY)
    );
    X_INV \IRDY/SRMUX (
      .I (N_RST),
      .O (\IRDY/SRNOT )
    );
    X_BUF \IRDY/IMUX (
      .I (\IRDY/IBUF ),
      .O (N_IRDY)
    );
    X_INV \IRDY/TRIMUX (
      .I (\bridge/out_bckp_frame_en_out ),
      .O (\IRDY/TNOT )
    );
    X_AND2 \IRDY/OUTBUF_GTS_AND_176 (
      .I0 (\IRDY/ENABLE ),
      .I1 (\IRDY/OUTBUF_GTS_AND_1_INV ),
      .O (\IRDY/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_irdy_reg_out_reg (
      .I (\IRDY/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\IRDY/IFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/in_reg_irdy_out )
    );
    X_OR2 \IRDY/IFF/ASYNC_FF_GSR_OR_177 (
      .I0 (\IRDY/SRNOT ),
      .I1 (GSR),
      .O (\IRDY/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/irdy_iob/dat_out_reg (
      .I (\bridge/pci_mux_irdy_in ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\IRDY/OFF/ASYNC_FF_GSR_OR ),
      .O (IRDY_out)
    );
    X_OR2 \IRDY/OFF/ASYNC_FF_GSR_OR_178 (
      .I0 (\IRDY/SRNOT ),
      .I1 (GSR),
      .O (\IRDY/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/irdy_iob/en_out_reg (
      .I (\IRDY/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\IRDY/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (IRDY_en)
    );
    X_OR2 \IRDY/TFF/ASYNC_FF_GSR_OR_179 (
      .I0 (\IRDY/SRNOT ),
      .I1 (GSR),
      .O (\IRDY/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<13>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[13]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<12> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [12]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [12])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<13> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [13]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [13])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[13]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<20>/DELAY (
      .I (N_AD[20]),
      .O (\AD[20]/IDELAY )
    );
    X_BUF \C15413/IBUF (
      .I (AD[20]),
      .O (N_AD[20])
    );
    X_INV \AD<20>/ENABLEINV (
      .I (AD_en[20]),
      .O (\AD[20]/ENABLE )
    );
    X_TRI \C15413/OBUFT (
      .I (AD_out[20]),
      .O (AD[20]),
      .CTL (\AD[20]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<20>/KEEPER (
      .O (\AD[20]/KEEPER )
    );
    X_BPAD \AD<20>/PAD (
      .PAD (AD[20])
    );
    X_INV \AD<20>/SRMUX (
      .I (N_RST),
      .O (\AD[20]/SRNOT )
    );
    X_BUF \AD<20>/OMUX (
      .I (\bridge/output_backup/C3/N126 ),
      .O (\AD[20]/OD )
    );
    X_AND2 \AD<20>/OUTBUF_GTS_AND (
      .I0 (\AD[20]/ENABLE ),
      .I1 (\AD[20]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[20]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<20> (
      .I (\AD[20]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[20]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [20])
    );
    X_OR2 \AD<20>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[20]/SRNOT ),
      .I1 (GSR),
      .O (\AD[20]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob20/dat_out_reg (
      .I (\AD[20]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mhigh ),
      .SET (GND),
      .RST (\AD[20]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[20])
    );
    X_OR2 \AD<20>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[20]/SRNOT ),
      .I1 (GSR),
      .O (\AD[20]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob20/en_out_reg (
      .I (N12330),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[20]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[20])
    );
    X_OR2 \AD<20>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[20]/SRNOT ),
      .I1 (GSR),
      .O (\AD[20]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \SERR/ENABLEINV (
      .I (SERR_en),
      .O (\SERR/ENABLE )
    );
    X_TRI C_SERR(
      .I (SERR_out),
      .O (SERR),
      .CTL (\SERR/OUTBUF_GTS_AND )
    );
    X_KEEPER \SERR/KEEPER_180 (
      .O (\SERR/KEEPER )
    );
    X_OPAD \SERR/PAD (
      .PAD (SERR)
    );
    X_INV \SERR/SRMUX (
      .I (N_RST),
      .O (\SERR/SRNOT )
    );
    X_BUF \SERR/OMUX (
      .I (N12029),
      .O (\SERR/OD )
    );
    X_INV \SERR/TRIMUX (
      .I (\bridge/pci_mux_serr_en_in ),
      .O (\SERR/TNOT )
    );
    X_AND2 \SERR/OUTBUF_GTS_AND_181 (
      .I0 (\SERR/ENABLE ),
      .I1 (\SERR/OUTBUF_GTS_AND_1_INV ),
      .O (\SERR/OUTBUF_GTS_AND )
    );
    X_FF \bridge/pci_io_mux/serr_iob/dat_out_reg (
      .I (\SERR/OD ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\SERR/OFF/ASYNC_FF_GSR_OR ),
      .O (SERR_out)
    );
    X_OR2 \SERR/OFF/ASYNC_FF_GSR_OR_182 (
      .I0 (\SERR/SRNOT ),
      .I1 (GSR),
      .O (\SERR/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/serr_iob/en_out_reg (
      .I (\SERR/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\SERR/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (SERR_en)
    );
    X_OR2 \SERR/TFF/ASYNC_FF_GSR_OR_183 (
      .I0 (\SERR/SRNOT ),
      .I1 (GSR),
      .O (\SERR/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<21>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[21]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<20> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [20]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[21]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [20])
    );
    X_OR2 \CRT/pix_start_addr<21>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[21]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[21]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<21> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [21]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[21]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [21])
    );
    X_OR2 \CRT/pix_start_addr<21>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[21]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[21]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<19>/DELAY (
      .I (N_AD[19]),
      .O (\AD[19]/IDELAY )
    );
    X_BUF \C15414/IBUF (
      .I (AD[19]),
      .O (N_AD[19])
    );
    X_INV \AD<19>/ENABLEINV (
      .I (AD_en[19]),
      .O (\AD[19]/ENABLE )
    );
    X_TRI \C15414/OBUFT (
      .I (AD_out[19]),
      .O (AD[19]),
      .CTL (\AD[19]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<19>/KEEPER (
      .O (\AD[19]/KEEPER )
    );
    X_BPAD \AD<19>/PAD (
      .PAD (AD[19])
    );
    X_INV \AD<19>/SRMUX (
      .I (N_RST),
      .O (\AD[19]/SRNOT )
    );
    X_BUF \AD<19>/OMUX (
      .I (\bridge/output_backup/C3/N120 ),
      .O (\AD[19]/OD )
    );
    X_AND2 \AD<19>/OUTBUF_GTS_AND (
      .I0 (\AD[19]/ENABLE ),
      .I1 (\AD[19]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[19]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<19> (
      .I (\AD[19]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[19]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [19])
    );
    X_OR2 \AD<19>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[19]/SRNOT ),
      .I1 (GSR),
      .O (\AD[19]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob19/dat_out_reg (
      .I (\AD[19]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mhigh ),
      .SET (GND),
      .RST (\AD[19]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[19])
    );
    X_OR2 \AD<19>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[19]/SRNOT ),
      .I1 (GSR),
      .O (\AD[19]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob19/en_out_reg (
      .I (N12330),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[19]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[19])
    );
    X_OR2 \AD<19>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[19]/SRNOT ),
      .I1 (GSR),
      .O (\AD[19]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<13>/DELAY (
      .I (N_AD[13]),
      .O (\AD[13]/IDELAY )
    );
    X_BUF \C15420/IBUF (
      .I (AD[13]),
      .O (N_AD[13])
    );
    X_INV \AD<13>/ENABLEINV (
      .I (AD_en[13]),
      .O (\AD[13]/ENABLE )
    );
    X_TRI \C15420/OBUFT (
      .I (AD_out[13]),
      .O (AD[13]),
      .CTL (\AD[13]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<13>/KEEPER (
      .O (\AD[13]/KEEPER )
    );
    X_BPAD \AD<13>/PAD (
      .PAD (AD[13])
    );
    X_INV \AD<13>/SRMUX (
      .I (N_RST),
      .O (\AD[13]/SRNOT )
    );
    X_BUF \AD<13>/OMUX (
      .I (\bridge/output_backup/C3/N84 ),
      .O (\AD[13]/OD )
    );
    X_AND2 \AD<13>/OUTBUF_GTS_AND (
      .I0 (\AD[13]/ENABLE ),
      .I1 (\AD[13]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[13]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<13> (
      .I (\AD[13]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[13]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [13])
    );
    X_OR2 \AD<13>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[13]/SRNOT ),
      .I1 (GSR),
      .O (\AD[13]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob13/dat_out_reg (
      .I (\AD[13]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mlow ),
      .SET (GND),
      .RST (\AD[13]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[13])
    );
    X_OR2 \AD<13>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[13]/SRNOT ),
      .I1 (GSR),
      .O (\AD[13]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob13/en_out_reg (
      .I (N12322),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[13]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[13])
    );
    X_OR2 \AD<13>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[13]/SRNOT ),
      .I1 (GSR),
      .O (\AD[13]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<13>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[13]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<12> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [12]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[13]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [12])
    );
    X_OR2 \CRT/pix_start_addr<13>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[13]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[13]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<13> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [13]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[13]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [13])
    );
    X_OR2 \CRT/pix_start_addr<13>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[13]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[13]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \C15451/IBUF (
      .I (PAR),
      .O (\PAR/IBUF )
    );
    X_INV \PAR/ENABLEINV (
      .I (PAR_en),
      .O (\PAR/ENABLE )
    );
    X_TRI \C15451/OBUFT (
      .I (PAR_out),
      .O (PAR),
      .CTL (\PAR/OUTBUF_GTS_AND )
    );
    X_KEEPER \PAR/KEEPER_184 (
      .O (\PAR/KEEPER )
    );
    X_BPAD \PAR/PAD (
      .PAD (PAR)
    );
    X_INV \PAR/SRMUX (
      .I (N_RST),
      .O (\PAR/SRNOT )
    );
    X_BUF \PAR/IMUX (
      .I (\PAR/IBUF ),
      .O (N_PAR)
    );
    X_INV \PAR/TRIMUX (
      .I (\bridge/pci_mux_par_en_in ),
      .O (\PAR/TNOT )
    );
    X_AND2 \PAR/OUTBUF_GTS_AND_185 (
      .I0 (\PAR/ENABLE ),
      .I1 (\PAR/OUTBUF_GTS_AND_1_INV ),
      .O (\PAR/OUTBUF_GTS_AND )
    );
    X_FF \bridge/pci_io_mux/par_iob/dat_out_reg (
      .I (\bridge/pci_mux_par_in ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\PAR/OFF/ASYNC_FF_GSR_OR ),
      .O (PAR_out)
    );
    X_OR2 \PAR/OFF/ASYNC_FF_GSR_OR_186 (
      .I0 (\PAR/SRNOT ),
      .I1 (GSR),
      .O (\PAR/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/par_iob/en_out_reg (
      .I (\PAR/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\PAR/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (PAR_en)
    );
    X_OR2 \PAR/TFF/ASYNC_FF_GSR_OR_187 (
      .I0 (\PAR/SRNOT ),
      .I1 (GSR),
      .O (\PAR/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<18>/DELAY (
      .I (N_AD[18]),
      .O (\AD[18]/IDELAY )
    );
    X_BUF \C15415/IBUF (
      .I (AD[18]),
      .O (N_AD[18])
    );
    X_INV \AD<18>/ENABLEINV (
      .I (AD_en[18]),
      .O (\AD[18]/ENABLE )
    );
    X_TRI \C15415/OBUFT (
      .I (AD_out[18]),
      .O (AD[18]),
      .CTL (\AD[18]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<18>/KEEPER (
      .O (\AD[18]/KEEPER )
    );
    X_BPAD \AD<18>/PAD (
      .PAD (AD[18])
    );
    X_INV \AD<18>/SRMUX (
      .I (N_RST),
      .O (\AD[18]/SRNOT )
    );
    X_BUF \AD<18>/OMUX (
      .I (\bridge/output_backup/C3/N114 ),
      .O (\AD[18]/OD )
    );
    X_AND2 \AD<18>/OUTBUF_GTS_AND (
      .I0 (\AD[18]/ENABLE ),
      .I1 (\AD[18]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[18]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<18> (
      .I (\AD[18]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[18]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [18])
    );
    X_OR2 \AD<18>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[18]/SRNOT ),
      .I1 (GSR),
      .O (\AD[18]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob18/dat_out_reg (
      .I (\AD[18]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mhigh ),
      .SET (GND),
      .RST (\AD[18]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[18])
    );
    X_OR2 \AD<18>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[18]/SRNOT ),
      .I1 (GSR),
      .O (\AD[18]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob18/en_out_reg (
      .I (N12330),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[18]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[18])
    );
    X_OR2 \AD<18>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[18]/SRNOT ),
      .I1 (GSR),
      .O (\AD[18]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<12>/DELAY (
      .I (N_AD[12]),
      .O (\AD[12]/IDELAY )
    );
    X_BUF \C15421/IBUF (
      .I (AD[12]),
      .O (N_AD[12])
    );
    X_INV \AD<12>/ENABLEINV (
      .I (AD_en[12]),
      .O (\AD[12]/ENABLE )
    );
    X_TRI \C15421/OBUFT (
      .I (AD_out[12]),
      .O (AD[12]),
      .CTL (\AD[12]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<12>/KEEPER (
      .O (\AD[12]/KEEPER )
    );
    X_BPAD \AD<12>/PAD (
      .PAD (AD[12])
    );
    X_INV \AD<12>/SRMUX (
      .I (N_RST),
      .O (\AD[12]/SRNOT )
    );
    X_BUF \AD<12>/OMUX (
      .I (\bridge/output_backup/C3/N78 ),
      .O (\AD[12]/OD )
    );
    X_AND2 \AD<12>/OUTBUF_GTS_AND (
      .I0 (\AD[12]/ENABLE ),
      .I1 (\AD[12]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[12]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<12> (
      .I (\AD[12]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[12]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [12])
    );
    X_OR2 \AD<12>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[12]/SRNOT ),
      .I1 (GSR),
      .O (\AD[12]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob12/dat_out_reg (
      .I (\AD[12]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mlow ),
      .SET (GND),
      .RST (\AD[12]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[12])
    );
    X_OR2 \AD<12>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[12]/SRNOT ),
      .I1 (GSR),
      .O (\AD[12]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob12/en_out_reg (
      .I (N12322),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[12]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[12])
    );
    X_OR2 \AD<12>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[12]/SRNOT ),
      .I1 (GSR),
      .O (\AD[12]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \CBE<1>/DELAY (
      .I (\CBE[1]/IBUF ),
      .O (\CBE[1]/IDELAY )
    );
    X_BUF \C15436/IBUF (
      .I (CBE[1]),
      .O (\CBE[1]/IBUF )
    );
    X_INV \CBE<1>/ENABLEINV (
      .I (CBE_en[1]),
      .O (\CBE[1]/ENABLE )
    );
    X_TRI \C15436/OBUFT (
      .I (CBE_out[1]),
      .O (CBE[1]),
      .CTL (\CBE[1]/OUTBUF_GTS_AND )
    );
    X_KEEPER \CBE<1>/KEEPER (
      .O (\CBE[1]/KEEPER )
    );
    X_BPAD \CBE<1>/PAD (
      .PAD (CBE[1])
    );
    X_INV \CBE<1>/SRMUX (
      .I (N_RST),
      .O (\CBE[1]/SRNOT )
    );
    X_BUF \CBE<1>/IMUX (
      .I (\CBE[1]/IBUF ),
      .O (N_CBE[1])
    );
    X_BUF \CBE<1>/OMUX (
      .I (\bridge/pci_mux_cbe_in [1]),
      .O (\CBE[1]/OD )
    );
    X_INV \CBE<1>/TRIMUX (
      .I (\bridge/pci_mux_cbe_en_in ),
      .O (\CBE[1]/TNOT )
    );
    X_AND2 \CBE<1>/OUTBUF_GTS_AND (
      .I0 (\CBE[1]/ENABLE ),
      .I1 (\CBE[1]/OUTBUF_GTS_AND_1_INV ),
      .O (\CBE[1]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_cbe_reg_out_reg<1> (
      .I (\CBE[1]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CBE[1]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/in_reg_cbe_out [1])
    );
    X_OR2 \CBE<1>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[1]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[1]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/cbe_iob1/dat_out_reg (
      .I (\CBE[1]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_mas_load_in ),
      .SET (GND),
      .RST (\CBE[1]/OFF/ASYNC_FF_GSR_OR ),
      .O (CBE_out[1])
    );
    X_OR2 \CBE<1>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[1]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[1]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/cbe_iob1/en_out_reg (
      .I (\CBE[1]/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\CBE[1]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (CBE_en[1])
    );
    X_OR2 \CBE<1>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[1]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[1]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \TRDY/DELAY (
      .I (\TRDY/IBUF ),
      .O (\TRDY/IDELAY )
    );
    X_BUF \C15449/IBUF (
      .I (TRDY),
      .O (\TRDY/IBUF )
    );
    X_INV \TRDY/ENABLEINV (
      .I (TRDY_en),
      .O (\TRDY/ENABLE )
    );
    X_TRI \C15449/OBUFT (
      .I (TRDY_out),
      .O (TRDY),
      .CTL (\TRDY/OUTBUF_GTS_AND )
    );
    X_KEEPER \TRDY/KEEPER_188 (
      .O (\TRDY/KEEPER )
    );
    X_BPAD \TRDY/PAD (
      .PAD (TRDY)
    );
    X_INV \TRDY/SRMUX (
      .I (N_RST),
      .O (\TRDY/SRNOT )
    );
    X_BUF \TRDY/IMUX (
      .I (\TRDY/IBUF ),
      .O (N_TRDY)
    );
    X_INV \TRDY/TRIMUX (
      .I (\bridge/pciu_pciif_devsel_en_out ),
      .O (\TRDY/TNOT )
    );
    X_AND2 \TRDY/OUTBUF_GTS_AND_189 (
      .I0 (\TRDY/ENABLE ),
      .I1 (\TRDY/OUTBUF_GTS_AND_1_INV ),
      .O (\TRDY/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_trdy_reg_out_reg (
      .I (\TRDY/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\TRDY/IFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/in_reg_trdy_out )
    );
    X_OR2 \TRDY/IFF/ASYNC_FF_GSR_OR_190 (
      .I0 (\TRDY/SRNOT ),
      .I1 (GSR),
      .O (\TRDY/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/trdy_iob/dat_out_reg (
      .I (N12472),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\TRDY/OFF/ASYNC_FF_GSR_OR ),
      .O (TRDY_out)
    );
    X_OR2 \TRDY/OFF/ASYNC_FF_GSR_OR_191 (
      .I0 (\TRDY/SRNOT ),
      .I1 (GSR),
      .O (\TRDY/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/trdy_iob/en_out_reg (
      .I (\TRDY/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\TRDY/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (TRDY_en)
    );
    X_OR2 \TRDY/TFF/ASYNC_FF_GSR_OR_192 (
      .I0 (\TRDY/SRNOT ),
      .I1 (GSR),
      .O (\TRDY/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<11>/DELAY (
      .I (N_AD[11]),
      .O (\AD[11]/IDELAY )
    );
    X_BUF \C15422/IBUF (
      .I (AD[11]),
      .O (N_AD[11])
    );
    X_INV \AD<11>/ENABLEINV (
      .I (AD_en[11]),
      .O (\AD[11]/ENABLE )
    );
    X_TRI \C15422/OBUFT (
      .I (AD_out[11]),
      .O (AD[11]),
      .CTL (\AD[11]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<11>/KEEPER (
      .O (\AD[11]/KEEPER )
    );
    X_BPAD \AD<11>/PAD (
      .PAD (AD[11])
    );
    X_INV \AD<11>/SRMUX (
      .I (N_RST),
      .O (\AD[11]/SRNOT )
    );
    X_BUF \AD<11>/OMUX (
      .I (\bridge/output_backup/C3/N72 ),
      .O (\AD[11]/OD )
    );
    X_AND2 \AD<11>/OUTBUF_GTS_AND (
      .I0 (\AD[11]/ENABLE ),
      .I1 (\AD[11]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[11]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<11> (
      .I (\AD[11]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[11]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [11])
    );
    X_OR2 \AD<11>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[11]/SRNOT ),
      .I1 (GSR),
      .O (\AD[11]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob11/dat_out_reg (
      .I (\AD[11]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mlow ),
      .SET (GND),
      .RST (\AD[11]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[11])
    );
    X_OR2 \AD<11>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[11]/SRNOT ),
      .I1 (GSR),
      .O (\AD[11]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob11/en_out_reg (
      .I (N12322),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[11]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[11])
    );
    X_OR2 \AD<11>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[11]/SRNOT ),
      .I1 (GSR),
      .O (\AD[11]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<15>/DELAY (
      .I (N_AD[15]),
      .O (\AD[15]/IDELAY )
    );
    X_BUF \C15418/IBUF (
      .I (AD[15]),
      .O (N_AD[15])
    );
    X_INV \AD<15>/ENABLEINV (
      .I (AD_en[15]),
      .O (\AD[15]/ENABLE )
    );
    X_TRI \C15418/OBUFT (
      .I (AD_out[15]),
      .O (AD[15]),
      .CTL (\AD[15]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<15>/KEEPER (
      .O (\AD[15]/KEEPER )
    );
    X_BPAD \AD<15>/PAD (
      .PAD (AD[15])
    );
    X_INV \AD<15>/SRMUX (
      .I (N_RST),
      .O (\AD[15]/SRNOT )
    );
    X_BUF \AD<15>/OMUX (
      .I (\bridge/output_backup/C3/N96 ),
      .O (\AD[15]/OD )
    );
    X_AND2 \AD<15>/OUTBUF_GTS_AND (
      .I0 (\AD[15]/ENABLE ),
      .I1 (\AD[15]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[15]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<15> (
      .I (\AD[15]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[15]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [15])
    );
    X_OR2 \AD<15>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[15]/SRNOT ),
      .I1 (GSR),
      .O (\AD[15]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob15/dat_out_reg (
      .I (\AD[15]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mlow ),
      .SET (GND),
      .RST (\AD[15]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[15])
    );
    X_OR2 \AD<15>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[15]/SRNOT ),
      .I1 (GSR),
      .O (\AD[15]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob15/en_out_reg (
      .I (N12322),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[15]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[15])
    );
    X_OR2 \AD<15>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[15]/SRNOT ),
      .I1 (GSR),
      .O (\AD[15]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<14>/DELAY (
      .I (N_AD[14]),
      .O (\AD[14]/IDELAY )
    );
    X_BUF \C15419/IBUF (
      .I (AD[14]),
      .O (N_AD[14])
    );
    X_INV \AD<14>/ENABLEINV (
      .I (AD_en[14]),
      .O (\AD[14]/ENABLE )
    );
    X_TRI \C15419/OBUFT (
      .I (AD_out[14]),
      .O (AD[14]),
      .CTL (\AD[14]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<14>/KEEPER (
      .O (\AD[14]/KEEPER )
    );
    X_BPAD \AD<14>/PAD (
      .PAD (AD[14])
    );
    X_INV \AD<14>/SRMUX (
      .I (N_RST),
      .O (\AD[14]/SRNOT )
    );
    X_BUF \AD<14>/OMUX (
      .I (\bridge/output_backup/C3/N90 ),
      .O (\AD[14]/OD )
    );
    X_AND2 \AD<14>/OUTBUF_GTS_AND (
      .I0 (\AD[14]/ENABLE ),
      .I1 (\AD[14]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[14]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<14> (
      .I (\AD[14]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[14]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [14])
    );
    X_OR2 \AD<14>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[14]/SRNOT ),
      .I1 (GSR),
      .O (\AD[14]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob14/dat_out_reg (
      .I (\AD[14]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mlow ),
      .SET (GND),
      .RST (\AD[14]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[14])
    );
    X_OR2 \AD<14>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[14]/SRNOT ),
      .I1 (GSR),
      .O (\AD[14]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob14/en_out_reg (
      .I (N12322),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[14]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[14])
    );
    X_OR2 \AD<14>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[14]/SRNOT ),
      .I1 (GSR),
      .O (\AD[14]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \DEVSEL/DELAY (
      .I (\DEVSEL/IBUF ),
      .O (\DEVSEL/IDELAY )
    );
    X_BUF \C15448/IBUF (
      .I (DEVSEL),
      .O (\DEVSEL/IBUF )
    );
    X_INV \DEVSEL/ENABLEINV (
      .I (DEVSEL_en),
      .O (\DEVSEL/ENABLE )
    );
    X_TRI \C15448/OBUFT (
      .I (DEVSEL_out),
      .O (DEVSEL),
      .CTL (\DEVSEL/OUTBUF_GTS_AND )
    );
    X_KEEPER \DEVSEL/KEEPER_193 (
      .O (\DEVSEL/KEEPER )
    );
    X_BPAD \DEVSEL/PAD (
      .PAD (DEVSEL)
    );
    X_INV \DEVSEL/SRMUX (
      .I (N_RST),
      .O (\DEVSEL/SRNOT )
    );
    X_BUF \DEVSEL/IMUX (
      .I (\DEVSEL/IBUF ),
      .O (N_DEVSEL)
    );
    X_INV \DEVSEL/TRIMUX (
      .I (\bridge/pciu_pciif_devsel_en_out ),
      .O (\DEVSEL/TNOT )
    );
    X_AND2 \DEVSEL/OUTBUF_GTS_AND_194 (
      .I0 (\DEVSEL/ENABLE ),
      .I1 (\DEVSEL/OUTBUF_GTS_AND_1_INV ),
      .O (\DEVSEL/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_devsel_reg_out_reg (
      .I (\DEVSEL/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\DEVSEL/IFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/in_reg_devsel_out )
    );
    X_OR2 \DEVSEL/IFF/ASYNC_FF_GSR_OR_195 (
      .I0 (\DEVSEL/SRNOT ),
      .I1 (GSR),
      .O (\DEVSEL/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/devsel_iob/dat_out_reg (
      .I (N12474),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\DEVSEL/OFF/ASYNC_FF_GSR_OR ),
      .O (DEVSEL_out)
    );
    X_OR2 \DEVSEL/OFF/ASYNC_FF_GSR_OR_196 (
      .I0 (\DEVSEL/SRNOT ),
      .I1 (GSR),
      .O (\DEVSEL/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/devsel_iob/en_out_reg (
      .I (\DEVSEL/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\DEVSEL/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (DEVSEL_en)
    );
    X_OR2 \DEVSEL/TFF/ASYNC_FF_GSR_OR_197 (
      .I0 (\DEVSEL/SRNOT ),
      .I1 (GSR),
      .O (\DEVSEL/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<10>/DELAY (
      .I (N_AD[10]),
      .O (\AD[10]/IDELAY )
    );
    X_BUF \C15423/IBUF (
      .I (AD[10]),
      .O (N_AD[10])
    );
    X_INV \AD<10>/ENABLEINV (
      .I (AD_en[10]),
      .O (\AD[10]/ENABLE )
    );
    X_TRI \C15423/OBUFT (
      .I (AD_out[10]),
      .O (AD[10]),
      .CTL (\AD[10]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<10>/KEEPER (
      .O (\AD[10]/KEEPER )
    );
    X_BPAD \AD<10>/PAD (
      .PAD (AD[10])
    );
    X_INV \AD<10>/SRMUX (
      .I (N_RST),
      .O (\AD[10]/SRNOT )
    );
    X_BUF \AD<10>/OMUX (
      .I (\bridge/output_backup/C3/N66 ),
      .O (\AD[10]/OD )
    );
    X_AND2 \AD<10>/OUTBUF_GTS_AND (
      .I0 (\AD[10]/ENABLE ),
      .I1 (\AD[10]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[10]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<10> (
      .I (\AD[10]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[10]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [10])
    );
    X_OR2 \AD<10>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[10]/SRNOT ),
      .I1 (GSR),
      .O (\AD[10]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob10/dat_out_reg (
      .I (\AD[10]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mlow ),
      .SET (GND),
      .RST (\AD[10]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[10])
    );
    X_OR2 \AD<10>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[10]/SRNOT ),
      .I1 (GSR),
      .O (\AD[10]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob10/en_out_reg (
      .I (N12322),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[10]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[10])
    );
    X_OR2 \AD<10>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[10]/SRNOT ),
      .I1 (GSR),
      .O (\AD[10]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<3>/DELAY (
      .I (N_AD[3]),
      .O (\AD[3]/IDELAY )
    );
    X_BUF \C15430/IBUF (
      .I (AD[3]),
      .O (N_AD[3])
    );
    X_INV \AD<3>/ENABLEINV (
      .I (AD_en[3]),
      .O (\AD[3]/ENABLE )
    );
    X_TRI \C15430/OBUFT (
      .I (AD_out[3]),
      .O (AD[3]),
      .CTL (\AD[3]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<3>/KEEPER (
      .O (\AD[3]/KEEPER )
    );
    X_BPAD \AD<3>/PAD (
      .PAD (AD[3])
    );
    X_INV \AD<3>/SRMUX (
      .I (N_RST),
      .O (\AD[3]/SRNOT )
    );
    X_BUF \AD<3>/OMUX (
      .I (\bridge/output_backup/C3/N24 ),
      .O (\AD[3]/OD )
    );
    X_AND2 \AD<3>/OUTBUF_GTS_AND (
      .I0 (\AD[3]/ENABLE ),
      .I1 (\AD[3]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[3]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<3> (
      .I (\AD[3]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[3]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [3])
    );
    X_OR2 \AD<3>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[3]/SRNOT ),
      .I1 (GSR),
      .O (\AD[3]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob3/dat_out_reg (
      .I (\AD[3]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_low ),
      .SET (GND),
      .RST (\AD[3]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[3])
    );
    X_OR2 \AD<3>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[3]/SRNOT ),
      .I1 (GSR),
      .O (\AD[3]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob3/en_out_reg (
      .I (N12314),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[3]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[3])
    );
    X_OR2 \AD<3>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[3]/SRNOT ),
      .I1 (GSR),
      .O (\AD[3]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<9>/DELAY (
      .I (N_AD[9]),
      .O (\AD[9]/IDELAY )
    );
    X_BUF \C15424/IBUF (
      .I (AD[9]),
      .O (N_AD[9])
    );
    X_INV \AD<9>/ENABLEINV (
      .I (AD_en[9]),
      .O (\AD[9]/ENABLE )
    );
    X_TRI \C15424/OBUFT (
      .I (AD_out[9]),
      .O (AD[9]),
      .CTL (\AD[9]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<9>/KEEPER (
      .O (\AD[9]/KEEPER )
    );
    X_BPAD \AD<9>/PAD (
      .PAD (AD[9])
    );
    X_INV \AD<9>/SRMUX (
      .I (N_RST),
      .O (\AD[9]/SRNOT )
    );
    X_BUF \AD<9>/OMUX (
      .I (\bridge/output_backup/C3/N60 ),
      .O (\AD[9]/OD )
    );
    X_AND2 \AD<9>/OUTBUF_GTS_AND (
      .I0 (\AD[9]/ENABLE ),
      .I1 (\AD[9]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[9]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<9> (
      .I (\AD[9]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[9]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [9])
    );
    X_OR2 \AD<9>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[9]/SRNOT ),
      .I1 (GSR),
      .O (\AD[9]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob9/dat_out_reg (
      .I (\AD[9]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mlow ),
      .SET (GND),
      .RST (\AD[9]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[9])
    );
    X_OR2 \AD<9>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[9]/SRNOT ),
      .I1 (GSR),
      .O (\AD[9]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob9/en_out_reg (
      .I (N12322),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[9]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[9])
    );
    X_OR2 \AD<9>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[9]/SRNOT ),
      .I1 (GSR),
      .O (\AD[9]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<2>/DELAY (
      .I (N_AD[2]),
      .O (\AD[2]/IDELAY )
    );
    X_BUF \C15431/IBUF (
      .I (AD[2]),
      .O (N_AD[2])
    );
    X_INV \AD<2>/ENABLEINV (
      .I (AD_en[2]),
      .O (\AD[2]/ENABLE )
    );
    X_TRI \C15431/OBUFT (
      .I (AD_out[2]),
      .O (AD[2]),
      .CTL (\AD[2]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<2>/KEEPER (
      .O (\AD[2]/KEEPER )
    );
    X_BPAD \AD<2>/PAD (
      .PAD (AD[2])
    );
    X_INV \AD<2>/SRMUX (
      .I (N_RST),
      .O (\AD[2]/SRNOT )
    );
    X_BUF \AD<2>/OMUX (
      .I (\bridge/output_backup/C3/N18 ),
      .O (\AD[2]/OD )
    );
    X_AND2 \AD<2>/OUTBUF_GTS_AND (
      .I0 (\AD[2]/ENABLE ),
      .I1 (\AD[2]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[2]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<2> (
      .I (\AD[2]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[2]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [2])
    );
    X_OR2 \AD<2>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[2]/SRNOT ),
      .I1 (GSR),
      .O (\AD[2]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob2/dat_out_reg (
      .I (\AD[2]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_low ),
      .SET (GND),
      .RST (\AD[2]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[2])
    );
    X_OR2 \AD<2>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[2]/SRNOT ),
      .I1 (GSR),
      .O (\AD[2]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob2/en_out_reg (
      .I (N12314),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[2]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[2])
    );
    X_OR2 \AD<2>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[2]/SRNOT ),
      .I1 (GSR),
      .O (\AD[2]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<8>/DELAY (
      .I (N_AD[8]),
      .O (\AD[8]/IDELAY )
    );
    X_BUF \C15425/IBUF (
      .I (AD[8]),
      .O (N_AD[8])
    );
    X_INV \AD<8>/ENABLEINV (
      .I (AD_en[8]),
      .O (\AD[8]/ENABLE )
    );
    X_TRI \C15425/OBUFT (
      .I (AD_out[8]),
      .O (AD[8]),
      .CTL (\AD[8]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<8>/KEEPER (
      .O (\AD[8]/KEEPER )
    );
    X_BPAD \AD<8>/PAD (
      .PAD (AD[8])
    );
    X_INV \AD<8>/SRMUX (
      .I (N_RST),
      .O (\AD[8]/SRNOT )
    );
    X_BUF \AD<8>/OMUX (
      .I (\bridge/output_backup/C3/N54 ),
      .O (\AD[8]/OD )
    );
    X_AND2 \AD<8>/OUTBUF_GTS_AND (
      .I0 (\AD[8]/ENABLE ),
      .I1 (\AD[8]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[8]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<8> (
      .I (\AD[8]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[8]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [8])
    );
    X_OR2 \AD<8>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[8]/SRNOT ),
      .I1 (GSR),
      .O (\AD[8]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob8/dat_out_reg (
      .I (\AD[8]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_mlow ),
      .SET (GND),
      .RST (\AD[8]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[8])
    );
    X_OR2 \AD<8>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[8]/SRNOT ),
      .I1 (GSR),
      .O (\AD[8]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob8/en_out_reg (
      .I (N12322),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[8]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[8])
    );
    X_OR2 \AD<8>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[8]/SRNOT ),
      .I1 (GSR),
      .O (\AD[8]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/del_sync_addr_out<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync_addr_out[29]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<28> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [28]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [28])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/del_sync/addr_out_reg<29> (
      .I (\bridge/pci_target_unit/pcit_if_addr_out [29]),
      .CLK (CLK_BUFGPed),
      .CE (N12545),
      .SET (GND),
      .RST (\bridge/pci_target_unit/del_sync_addr_out[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync_addr_out [29])
    );
    X_OR2 \bridge/pci_target_unit/del_sync_addr_out<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/del_sync_addr_out[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/del_sync_addr_out[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<1>/DELAY (
      .I (N_AD[1]),
      .O (\AD[1]/IDELAY )
    );
    X_BUF \C15432/IBUF (
      .I (AD[1]),
      .O (N_AD[1])
    );
    X_INV \AD<1>/ENABLEINV (
      .I (AD_en[1]),
      .O (\AD[1]/ENABLE )
    );
    X_TRI \C15432/OBUFT (
      .I (AD_out[1]),
      .O (AD[1]),
      .CTL (\AD[1]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<1>/KEEPER (
      .O (\AD[1]/KEEPER )
    );
    X_BPAD \AD<1>/PAD (
      .PAD (AD[1])
    );
    X_INV \AD<1>/SRMUX (
      .I (N_RST),
      .O (\AD[1]/SRNOT )
    );
    X_AND2 \AD<1>/OUTBUF_GTS_AND (
      .I0 (\AD[1]/ENABLE ),
      .I1 (\AD[1]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[1]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<1> (
      .I (\AD[1]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[1]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [1])
    );
    X_OR2 \AD<1>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[1]/SRNOT ),
      .I1 (GSR),
      .O (\AD[1]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob1/dat_out_reg (
      .I (\bridge/output_backup/C3/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_low ),
      .SET (GND),
      .RST (\AD[1]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[1])
    );
    X_OR2 \AD<1>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[1]/SRNOT ),
      .I1 (GSR),
      .O (\AD[1]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob1/en_out_reg (
      .I (N12314),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[1]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[1])
    );
    X_OR2 \AD<1>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[1]/SRNOT ),
      .I1 (GSR),
      .O (\AD[1]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \CBE<0>/DELAY (
      .I (\CBE[0]/IBUF ),
      .O (\CBE[0]/IDELAY )
    );
    X_BUF \C15437/IBUF (
      .I (CBE[0]),
      .O (\CBE[0]/IBUF )
    );
    X_INV \CBE<0>/ENABLEINV (
      .I (CBE_en[0]),
      .O (\CBE[0]/ENABLE )
    );
    X_TRI \C15437/OBUFT (
      .I (CBE_out[0]),
      .O (CBE[0]),
      .CTL (\CBE[0]/OUTBUF_GTS_AND )
    );
    X_KEEPER \CBE<0>/KEEPER (
      .O (\CBE[0]/KEEPER )
    );
    X_BPAD \CBE<0>/PAD (
      .PAD (CBE[0])
    );
    X_INV \CBE<0>/SRMUX (
      .I (N_RST),
      .O (\CBE[0]/SRNOT )
    );
    X_BUF \CBE<0>/IMUX (
      .I (\CBE[0]/IBUF ),
      .O (N_CBE[0])
    );
    X_BUF \CBE<0>/OMUX (
      .I (\bridge/pci_mux_cbe_in [0]),
      .O (\CBE[0]/OD )
    );
    X_INV \CBE<0>/TRIMUX (
      .I (\bridge/pci_mux_cbe_en_in ),
      .O (\CBE[0]/TNOT )
    );
    X_AND2 \CBE<0>/OUTBUF_GTS_AND (
      .I0 (\CBE[0]/ENABLE ),
      .I1 (\CBE[0]/OUTBUF_GTS_AND_1_INV ),
      .O (\CBE[0]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_cbe_reg_out_reg<0> (
      .I (\CBE[0]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\CBE[0]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/in_reg_cbe_out [0])
    );
    X_OR2 \CBE<0>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[0]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[0]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/cbe_iob0/dat_out_reg (
      .I (\CBE[0]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_mux_mas_load_in ),
      .SET (GND),
      .RST (\CBE[0]/OFF/ASYNC_FF_GSR_OR ),
      .O (CBE_out[0])
    );
    X_OR2 \CBE<0>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[0]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[0]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/cbe_iob0/en_out_reg (
      .I (\CBE[0]/TNOT ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\CBE[0]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (CBE_en[0])
    );
    X_OR2 \CBE<0>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\CBE[0]/SRNOT ),
      .I1 (GSR),
      .O (\CBE[0]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<31>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[31]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<30> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [30]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [30])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<31> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [31]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [31])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[31]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<6>/DELAY (
      .I (N_AD[6]),
      .O (\AD[6]/IDELAY )
    );
    X_BUF \C15427/IBUF (
      .I (AD[6]),
      .O (N_AD[6])
    );
    X_INV \AD<6>/ENABLEINV (
      .I (AD_en[6]),
      .O (\AD[6]/ENABLE )
    );
    X_TRI \C15427/OBUFT (
      .I (AD_out[6]),
      .O (AD[6]),
      .CTL (\AD[6]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<6>/KEEPER (
      .O (\AD[6]/KEEPER )
    );
    X_BPAD \AD<6>/PAD (
      .PAD (AD[6])
    );
    X_INV \AD<6>/SRMUX (
      .I (N_RST),
      .O (\AD[6]/SRNOT )
    );
    X_BUF \AD<6>/OMUX (
      .I (\bridge/output_backup/C3/N42 ),
      .O (\AD[6]/OD )
    );
    X_AND2 \AD<6>/OUTBUF_GTS_AND (
      .I0 (\AD[6]/ENABLE ),
      .I1 (\AD[6]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[6]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<6> (
      .I (\AD[6]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[6]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [6])
    );
    X_OR2 \AD<6>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[6]/SRNOT ),
      .I1 (GSR),
      .O (\AD[6]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob6/dat_out_reg (
      .I (\AD[6]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_low ),
      .SET (GND),
      .RST (\AD[6]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[6])
    );
    X_OR2 \AD<6>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[6]/SRNOT ),
      .I1 (GSR),
      .O (\AD[6]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob6/en_out_reg (
      .I (N12314),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[6]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[6])
    );
    X_OR2 \AD<6>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[6]/SRNOT ),
      .I1 (GSR),
      .O (\AD[6]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<7>/DELAY (
      .I (N_AD[7]),
      .O (\AD[7]/IDELAY )
    );
    X_BUF \C15426/IBUF (
      .I (AD[7]),
      .O (N_AD[7])
    );
    X_INV \AD<7>/ENABLEINV (
      .I (AD_en[7]),
      .O (\AD[7]/ENABLE )
    );
    X_TRI \C15426/OBUFT (
      .I (AD_out[7]),
      .O (AD[7]),
      .CTL (\AD[7]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<7>/KEEPER (
      .O (\AD[7]/KEEPER )
    );
    X_BPAD \AD<7>/PAD (
      .PAD (AD[7])
    );
    X_INV \AD<7>/SRMUX (
      .I (N_RST),
      .O (\AD[7]/SRNOT )
    );
    X_BUF \AD<7>/OMUX (
      .I (\bridge/output_backup/C3/N48 ),
      .O (\AD[7]/OD )
    );
    X_AND2 \AD<7>/OUTBUF_GTS_AND (
      .I0 (\AD[7]/ENABLE ),
      .I1 (\AD[7]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[7]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<7> (
      .I (\AD[7]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[7]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [7])
    );
    X_OR2 \AD<7>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[7]/SRNOT ),
      .I1 (GSR),
      .O (\AD[7]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob7/dat_out_reg (
      .I (\AD[7]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_low ),
      .SET (GND),
      .RST (\AD[7]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[7])
    );
    X_OR2 \AD<7>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[7]/SRNOT ),
      .I1 (GSR),
      .O (\AD[7]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob7/en_out_reg (
      .I (N12314),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[7]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[7])
    );
    X_OR2 \AD<7>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[7]/SRNOT ),
      .I1 (GSR),
      .O (\AD[7]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<23>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[23]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<22> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [22]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [22])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<23> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [23]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [23])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[23]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<5>/DELAY (
      .I (N_AD[5]),
      .O (\AD[5]/IDELAY )
    );
    X_BUF \C15428/IBUF (
      .I (AD[5]),
      .O (N_AD[5])
    );
    X_INV \AD<5>/ENABLEINV (
      .I (AD_en[5]),
      .O (\AD[5]/ENABLE )
    );
    X_TRI \C15428/OBUFT (
      .I (AD_out[5]),
      .O (AD[5]),
      .CTL (\AD[5]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<5>/KEEPER (
      .O (\AD[5]/KEEPER )
    );
    X_BPAD \AD<5>/PAD (
      .PAD (AD[5])
    );
    X_INV \AD<5>/SRMUX (
      .I (N_RST),
      .O (\AD[5]/SRNOT )
    );
    X_BUF \AD<5>/OMUX (
      .I (\bridge/output_backup/C3/N36 ),
      .O (\AD[5]/OD )
    );
    X_AND2 \AD<5>/OUTBUF_GTS_AND (
      .I0 (\AD[5]/ENABLE ),
      .I1 (\AD[5]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[5]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<5> (
      .I (\AD[5]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[5]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [5])
    );
    X_OR2 \AD<5>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[5]/SRNOT ),
      .I1 (GSR),
      .O (\AD[5]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob5/dat_out_reg (
      .I (\AD[5]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_low ),
      .SET (GND),
      .RST (\AD[5]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[5])
    );
    X_OR2 \AD<5>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[5]/SRNOT ),
      .I1 (GSR),
      .O (\AD[5]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob5/en_out_reg (
      .I (N12314),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[5]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[5])
    );
    X_OR2 \AD<5>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[5]/SRNOT ),
      .I1 (GSR),
      .O (\AD[5]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF C_GNT(
      .I (GNT),
      .O (\GNT/IBUF )
    );
    X_KEEPER \GNT/KEEPER_198 (
      .O (\GNT/KEEPER )
    );
    X_IPAD \GNT/PAD (
      .PAD (GNT)
    );
    X_BUF \GNT/IMUX (
      .I (\GNT/IBUF ),
      .O (N_GNT)
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<15>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[15]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<14> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [14]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [14])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<15> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [15]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [15])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[15]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \HSYNC/KEEPER_199 (
      .O (\HSYNC/KEEPER )
    );
    X_OPAD \HSYNC/PAD (
      .PAD (HSYNC)
    );
    X_INV \HSYNC/SRMUX (
      .I (N_RST),
      .O (\HSYNC/SRNOT )
    );
    X_BUF \HSYNC/OMUX (
      .I (crt_hsync),
      .O (\HSYNC/OD )
    );
    X_BUF C_HSYNC(
      .I (N_HSYNC),
      .O (\HSYNC/OUTBUF_GTS_TRI )
    );
    X_TRI C_HSYNC_200(
      .I (\HSYNC/OUTBUF_GTS_TRI ),
      .O (HSYNC),
      .CTL (C_HSYNC_2_INV)
    );
    X_FF \crt_out_reg/hsync_out_reg (
      .I (\HSYNC/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\HSYNC/OFF/ASYNC_FF_GSR_OR ),
      .O (N_HSYNC)
    );
    X_OR2 \HSYNC/OFF/ASYNC_FF_GSR_OR_201 (
      .I0 (\HSYNC/SRNOT ),
      .I1 (GSR),
      .O (\HSYNC/OFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<4>/DELAY (
      .I (N_AD[4]),
      .O (\AD[4]/IDELAY )
    );
    X_BUF \C15429/IBUF (
      .I (AD[4]),
      .O (N_AD[4])
    );
    X_INV \AD<4>/ENABLEINV (
      .I (AD_en[4]),
      .O (\AD[4]/ENABLE )
    );
    X_TRI \C15429/OBUFT (
      .I (AD_out[4]),
      .O (AD[4]),
      .CTL (\AD[4]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<4>/KEEPER (
      .O (\AD[4]/KEEPER )
    );
    X_BPAD \AD<4>/PAD (
      .PAD (AD[4])
    );
    X_INV \AD<4>/SRMUX (
      .I (N_RST),
      .O (\AD[4]/SRNOT )
    );
    X_BUF \AD<4>/OMUX (
      .I (\bridge/output_backup/C3/N30 ),
      .O (\AD[4]/OD )
    );
    X_AND2 \AD<4>/OUTBUF_GTS_AND (
      .I0 (\AD[4]/ENABLE ),
      .I1 (\AD[4]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[4]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<4> (
      .I (\AD[4]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[4]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [4])
    );
    X_OR2 \AD<4>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[4]/SRNOT ),
      .I1 (GSR),
      .O (\AD[4]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob4/dat_out_reg (
      .I (\AD[4]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_low ),
      .SET (GND),
      .RST (\AD[4]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[4])
    );
    X_OR2 \AD<4>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[4]/SRNOT ),
      .I1 (GSR),
      .O (\AD[4]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob4/en_out_reg (
      .I (N12314),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[4]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[4])
    );
    X_OR2 \AD<4>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[4]/SRNOT ),
      .I1 (GSR),
      .O (\AD[4]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<31>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[31]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<30> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [30]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[31]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [30])
    );
    X_OR2 \CRT/pix_start_addr<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[31]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[31]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<31> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [31]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[31]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [31])
    );
    X_OR2 \CRT/pix_start_addr<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[31]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[31]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \REQ/ENABLEINV (
      .I (REQ_en),
      .O (\REQ/ENABLE )
    );
    X_TRI C_REQ(
      .I (REQ_out),
      .O (REQ),
      .CTL (\REQ/OUTBUF_GTS_AND )
    );
    X_KEEPER \REQ/KEEPER_202 (
      .O (\REQ/KEEPER )
    );
    X_OPAD \REQ/PAD (
      .PAD (REQ)
    );
    X_INV \REQ/SRMUX (
      .I (N_RST),
      .O (\REQ/SRNOT )
    );
    X_BUF \REQ/OMUX (
      .I (N12587),
      .O (\REQ/OD )
    );
    X_ZERO \REQ/LOGIC_ZERO_203 (
      .O (\REQ/LOGIC_ZERO )
    );
    X_AND2 \REQ/OUTBUF_GTS_AND_204 (
      .I0 (\REQ/ENABLE ),
      .I1 (\REQ/OUTBUF_GTS_AND_1_INV ),
      .O (\REQ/OUTBUF_GTS_AND )
    );
    X_FF \bridge/pci_io_mux/req_iob/dat_out_reg (
      .I (\REQ/OD ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\REQ/OFF/ASYNC_FF_GSR_OR ),
      .O (REQ_out)
    );
    X_OR2 \REQ/OFF/ASYNC_FF_GSR_OR_205 (
      .I0 (\REQ/SRNOT ),
      .I1 (GSR),
      .O (\REQ/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/req_iob/en_out_reg (
      .I (\REQ/LOGIC_ZERO ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\REQ/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (REQ_en)
    );
    X_OR2 \REQ/TFF/ASYNC_FF_GSR_OR_206 (
      .I0 (\REQ/SRNOT ),
      .I1 (GSR),
      .O (\REQ/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<0>/DELAY (
      .I (N_AD[0]),
      .O (\AD[0]/IDELAY )
    );
    X_BUF \C15433/IBUF (
      .I (AD[0]),
      .O (N_AD[0])
    );
    X_INV \AD<0>/ENABLEINV (
      .I (AD_en[0]),
      .O (\AD[0]/ENABLE )
    );
    X_TRI \C15433/OBUFT (
      .I (AD_out[0]),
      .O (AD[0]),
      .CTL (\AD[0]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<0>/KEEPER (
      .O (\AD[0]/KEEPER )
    );
    X_BPAD \AD<0>/PAD (
      .PAD (AD[0])
    );
    X_INV \AD<0>/SRMUX (
      .I (N_RST),
      .O (\AD[0]/SRNOT )
    );
    X_BUF \AD<0>/OMUX (
      .I (\bridge/output_backup/C3/N6 ),
      .O (\AD[0]/OD )
    );
    X_AND2 \AD<0>/OUTBUF_GTS_AND (
      .I0 (\AD[0]/ENABLE ),
      .I1 (\AD[0]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[0]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<0> (
      .I (\AD[0]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[0]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [0])
    );
    X_OR2 \AD<0>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[0]/SRNOT ),
      .I1 (GSR),
      .O (\AD[0]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob0/dat_out_reg (
      .I (\AD[0]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_low ),
      .SET (GND),
      .RST (\AD[0]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[0])
    );
    X_OR2 \AD<0>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[0]/SRNOT ),
      .I1 (GSR),
      .O (\AD[0]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob0/en_out_reg (
      .I (N12314),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[0]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[0])
    );
    X_OR2 \AD<0>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[0]/SRNOT ),
      .I1 (GSR),
      .O (\AD[0]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<23>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[23]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<22> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [22]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[23]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [22])
    );
    X_OR2 \CRT/pix_start_addr<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[23]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[23]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<23> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [23]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[23]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [23])
    );
    X_OR2 \CRT/pix_start_addr<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[23]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[23]/FFX/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \VSYNC/KEEPER_207 (
      .O (\VSYNC/KEEPER )
    );
    X_OPAD \VSYNC/PAD (
      .PAD (VSYNC)
    );
    X_INV \VSYNC/SRMUX (
      .I (N_RST),
      .O (\VSYNC/SRNOT )
    );
    X_BUF \VSYNC/OMUX (
      .I (crt_vsync),
      .O (\VSYNC/OD )
    );
    X_BUF C_VSYNC(
      .I (N_VSYNC),
      .O (\VSYNC/OUTBUF_GTS_TRI )
    );
    X_TRI C_VSYNC_208(
      .I (\VSYNC/OUTBUF_GTS_TRI ),
      .O (VSYNC),
      .CTL (C_VSYNC_2_INV)
    );
    X_FF \crt_out_reg/vsync_out_reg (
      .I (\VSYNC/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\VSYNC/OFF/ASYNC_FF_GSR_OR ),
      .O (N_VSYNC)
    );
    X_OR2 \VSYNC/OFF/ASYNC_FF_GSR_OR_209 (
      .I0 (\VSYNC/SRNOT ),
      .I1 (GSR),
      .O (\VSYNC/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \LED/KEEPER_210 (
      .O (\LED/KEEPER )
    );
    X_OPAD \LED/PAD (
      .PAD (LED)
    );
    X_BUF \LED/OMUX (
      .I (N_LED),
      .O (\LED/OD )
    );
    X_BUF C_LED(
      .I (\LED/OD ),
      .O (\LED/OUTBUF_GTS_TRI )
    );
    X_TRI C_LED_211(
      .I (\LED/OUTBUF_GTS_TRI ),
      .O (LED),
      .CTL (C_LED_2_INV)
    );
    X_INV \CRT/pix_start_addr<15>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[15]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<14> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [14]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[15]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [14])
    );
    X_OR2 \CRT/pix_start_addr<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[15]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[15]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<15> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [15]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[15]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [15])
    );
    X_OR2 \CRT/pix_start_addr<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[15]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[15]/FFX/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<31>/DELAY (
      .I (N_AD[31]),
      .O (\AD[31]/IDELAY )
    );
    X_BUF \C15402/IBUF (
      .I (AD[31]),
      .O (N_AD[31])
    );
    X_INV \AD<31>/ENABLEINV (
      .I (AD_en[31]),
      .O (\AD[31]/ENABLE )
    );
    X_TRI \C15402/OBUFT (
      .I (AD_out[31]),
      .O (AD[31]),
      .CTL (\AD[31]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<31>/KEEPER (
      .O (\AD[31]/KEEPER )
    );
    X_BPAD \AD<31>/PAD (
      .PAD (AD[31])
    );
    X_INV \AD<31>/SRMUX (
      .I (N_RST),
      .O (\AD[31]/SRNOT )
    );
    X_AND2 \AD<31>/OUTBUF_GTS_AND (
      .I0 (\AD[31]/ENABLE ),
      .I1 (\AD[31]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[31]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<31> (
      .I (\AD[31]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[31]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [31])
    );
    X_OR2 \AD<31>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[31]/SRNOT ),
      .I1 (GSR),
      .O (\AD[31]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob31/dat_out_reg (
      .I (\bridge/output_backup/C3/N192 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_high ),
      .SET (GND),
      .RST (\AD[31]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[31])
    );
    X_OR2 \AD<31>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[31]/SRNOT ),
      .I1 (GSR),
      .O (\AD[31]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob31/en_out_reg (
      .I (N12338),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[31]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[31])
    );
    X_OR2 \AD<31>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[31]/SRNOT ),
      .I1 (GSR),
      .O (\AD[31]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<30>/DELAY (
      .I (N_AD[30]),
      .O (\AD[30]/IDELAY )
    );
    X_BUF \C15403/IBUF (
      .I (AD[30]),
      .O (N_AD[30])
    );
    X_INV \AD<30>/ENABLEINV (
      .I (AD_en[30]),
      .O (\AD[30]/ENABLE )
    );
    X_TRI \C15403/OBUFT (
      .I (AD_out[30]),
      .O (AD[30]),
      .CTL (\AD[30]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<30>/KEEPER (
      .O (\AD[30]/KEEPER )
    );
    X_BPAD \AD<30>/PAD (
      .PAD (AD[30])
    );
    X_INV \AD<30>/SRMUX (
      .I (N_RST),
      .O (\AD[30]/SRNOT )
    );
    X_AND2 \AD<30>/OUTBUF_GTS_AND (
      .I0 (\AD[30]/ENABLE ),
      .I1 (\AD[30]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[30]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<30> (
      .I (\AD[30]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[30]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [30])
    );
    X_OR2 \AD<30>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[30]/SRNOT ),
      .I1 (GSR),
      .O (\AD[30]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob30/dat_out_reg (
      .I (\bridge/output_backup/C3/N186 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_high ),
      .SET (GND),
      .RST (\AD[30]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[30])
    );
    X_OR2 \AD<30>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[30]/SRNOT ),
      .I1 (GSR),
      .O (\AD[30]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob30/en_out_reg (
      .I (N12338),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[30]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[30])
    );
    X_OR2 \AD<30>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[30]/SRNOT ),
      .I1 (GSR),
      .O (\AD[30]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<29>/DELAY (
      .I (N_AD[29]),
      .O (\AD[29]/IDELAY )
    );
    X_BUF \C15404/IBUF (
      .I (AD[29]),
      .O (N_AD[29])
    );
    X_INV \AD<29>/ENABLEINV (
      .I (AD_en[29]),
      .O (\AD[29]/ENABLE )
    );
    X_TRI \C15404/OBUFT (
      .I (AD_out[29]),
      .O (AD[29]),
      .CTL (\AD[29]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<29>/KEEPER (
      .O (\AD[29]/KEEPER )
    );
    X_BPAD \AD<29>/PAD (
      .PAD (AD[29])
    );
    X_INV \AD<29>/SRMUX (
      .I (N_RST),
      .O (\AD[29]/SRNOT )
    );
    X_BUF \AD<29>/OMUX (
      .I (\bridge/output_backup/C3/N180 ),
      .O (\AD[29]/OD )
    );
    X_AND2 \AD<29>/OUTBUF_GTS_AND (
      .I0 (\AD[29]/ENABLE ),
      .I1 (\AD[29]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[29]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<29> (
      .I (\AD[29]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[29]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [29])
    );
    X_OR2 \AD<29>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[29]/SRNOT ),
      .I1 (GSR),
      .O (\AD[29]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob29/dat_out_reg (
      .I (\AD[29]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_high ),
      .SET (GND),
      .RST (\AD[29]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[29])
    );
    X_OR2 \AD<29>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[29]/SRNOT ),
      .I1 (GSR),
      .O (\AD[29]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob29/en_out_reg (
      .I (N12338),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[29]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[29])
    );
    X_OR2 \AD<29>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[29]/SRNOT ),
      .I1 (GSR),
      .O (\AD[29]/TFF/ASYNC_FF_GSR_OR )
    );
    X_BUF \AD<28>/DELAY (
      .I (N_AD[28]),
      .O (\AD[28]/IDELAY )
    );
    X_BUF \C15405/IBUF (
      .I (AD[28]),
      .O (N_AD[28])
    );
    X_INV \AD<28>/ENABLEINV (
      .I (AD_en[28]),
      .O (\AD[28]/ENABLE )
    );
    X_TRI \C15405/OBUFT (
      .I (AD_out[28]),
      .O (AD[28]),
      .CTL (\AD[28]/OUTBUF_GTS_AND )
    );
    X_KEEPER \AD<28>/KEEPER (
      .O (\AD[28]/KEEPER )
    );
    X_BPAD \AD<28>/PAD (
      .PAD (AD[28])
    );
    X_INV \AD<28>/SRMUX (
      .I (N_RST),
      .O (\AD[28]/SRNOT )
    );
    X_BUF \AD<28>/OMUX (
      .I (\bridge/output_backup/C3/N174 ),
      .O (\AD[28]/OD )
    );
    X_AND2 \AD<28>/OUTBUF_GTS_AND (
      .I0 (\AD[28]/ENABLE ),
      .I1 (\AD[28]/OUTBUF_GTS_AND_1_INV ),
      .O (\AD[28]/OUTBUF_GTS_AND )
    );
    X_FF \bridge/input_register/pci_ad_reg_out_reg<28> (
      .I (\AD[28]/IDELAY ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\AD[28]/IFF/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/address1_in [28])
    );
    X_OR2 \AD<28>/IFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[28]/SRNOT ),
      .I1 (GSR),
      .O (\AD[28]/IFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob28/dat_out_reg (
      .I (\AD[28]/OD ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_io_mux/ad_load_ctrl_high ),
      .SET (GND),
      .RST (\AD[28]/OFF/ASYNC_FF_GSR_OR ),
      .O (AD_out[28])
    );
    X_OR2 \AD<28>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[28]/SRNOT ),
      .I1 (GSR),
      .O (\AD[28]/OFF/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_io_mux/ad_iob28/en_out_reg (
      .I (N12338),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (\AD[28]/TFF/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (AD_en[28])
    );
    X_OR2 \AD<28>/TFF/ASYNC_FF_GSR_OR (
      .I0 (\AD[28]/SRNOT ),
      .I1 (GSR),
      .O (\AD[28]/TFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_if_bc_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_bc_out[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_bc_reg<0> (
      .I (\bridge/in_reg_cbe_out [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_bc_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_bc_out [0])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_bc_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_bc_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_bc_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_bc_reg<1> (
      .I (\bridge/in_reg_cbe_out [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_bc_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_bc_out [1])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_bc_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_bc_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_bc_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<14>/KEEPER (
      .O (\RGB[14]/KEEPER )
    );
    X_OPAD \RGB<14>/PAD (
      .PAD (RGB[14])
    );
    X_INV \RGB<14>/SRMUX (
      .I (N_RST),
      .O (\RGB[14]/SRNOT )
    );
    X_BUF \RGB<14>/OMUX (
      .I (rgb_int[14]),
      .O (\RGB[14]/OD )
    );
    X_BUF \C_RGB<14> (
      .I (N_RGB[14]),
      .O (\RGB[14]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<14>_212 (
      .I (\RGB[14]/OUTBUF_GTS_TRI ),
      .O (RGB[14]),
      .CTL (\C_RGB[14]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<14> (
      .I (\RGB[14]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[14]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[14])
    );
    X_OR2 \RGB<14>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[14]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[14]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<7>/KEEPER (
      .O (\RGB[7]/KEEPER )
    );
    X_OPAD \RGB<7>/PAD (
      .PAD (RGB[7])
    );
    X_INV \RGB<7>/SRMUX (
      .I (N_RST),
      .O (\RGB[7]/SRNOT )
    );
    X_BUF \C_RGB<7> (
      .I (N_RGB[7]),
      .O (\RGB[7]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<7>_213 (
      .I (\RGB[7]/OUTBUF_GTS_TRI ),
      .O (RGB[7]),
      .CTL (\C_RGB[7]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<7> (
      .I (rgb_int[7]),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[7]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[7])
    );
    X_OR2 \RGB<7>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[7]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[7]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<15>/KEEPER (
      .O (\RGB[15]/KEEPER )
    );
    X_OPAD \RGB<15>/PAD (
      .PAD (RGB[15])
    );
    X_INV \RGB<15>/SRMUX (
      .I (N_RST),
      .O (\RGB[15]/SRNOT )
    );
    X_BUF \RGB<15>/OMUX (
      .I (rgb_int[15]),
      .O (\RGB[15]/OD )
    );
    X_BUF \C_RGB<15> (
      .I (N_RGB[15]),
      .O (\RGB[15]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<15>_214 (
      .I (\RGB[15]/OUTBUF_GTS_TRI ),
      .O (RGB[15]),
      .CTL (\C_RGB[15]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<15> (
      .I (\RGB[15]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[15]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[15])
    );
    X_OR2 \RGB<15>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[15]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[15]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<8>/KEEPER (
      .O (\RGB[8]/KEEPER )
    );
    X_OPAD \RGB<8>/PAD (
      .PAD (RGB[8])
    );
    X_INV \RGB<8>/SRMUX (
      .I (N_RST),
      .O (\RGB[8]/SRNOT )
    );
    X_BUF \RGB<8>/OMUX (
      .I (rgb_int[8]),
      .O (\RGB[8]/OD )
    );
    X_BUF \C_RGB<8> (
      .I (N_RGB[8]),
      .O (\RGB[8]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<8>_215 (
      .I (\RGB[8]/OUTBUF_GTS_TRI ),
      .O (RGB[8]),
      .CTL (\C_RGB[8]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<8> (
      .I (\RGB[8]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[8]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[8])
    );
    X_OR2 \RGB<8>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[8]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[8]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<9>/KEEPER (
      .O (\RGB[9]/KEEPER )
    );
    X_OPAD \RGB<9>/PAD (
      .PAD (RGB[9])
    );
    X_INV \RGB<9>/SRMUX (
      .I (N_RST),
      .O (\RGB[9]/SRNOT )
    );
    X_BUF \RGB<9>/OMUX (
      .I (rgb_int[9]),
      .O (\RGB[9]/OD )
    );
    X_BUF \C_RGB<9> (
      .I (N_RGB[9]),
      .O (\RGB[9]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<9>_216 (
      .I (\RGB[9]/OUTBUF_GTS_TRI ),
      .O (RGB[9]),
      .CTL (\C_RGB[9]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<9> (
      .I (\RGB[9]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[9]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[9])
    );
    X_OR2 \RGB<9>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[9]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[9]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<4>/KEEPER (
      .O (\RGB[4]/KEEPER )
    );
    X_OPAD \RGB<4>/PAD (
      .PAD (RGB[4])
    );
    X_INV \RGB<4>/SRMUX (
      .I (N_RST),
      .O (\RGB[4]/SRNOT )
    );
    X_BUF \RGB<4>/OMUX (
      .I (rgb_int[4]),
      .O (\RGB[4]/OD )
    );
    X_BUF \C_RGB<4> (
      .I (N_RGB[4]),
      .O (\RGB[4]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<4>_217 (
      .I (\RGB[4]/OUTBUF_GTS_TRI ),
      .O (RGB[4]),
      .CTL (\C_RGB[4]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<4> (
      .I (\RGB[4]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[4]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[4])
    );
    X_OR2 \RGB<4>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[4]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[4]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<5>/KEEPER (
      .O (\RGB[5]/KEEPER )
    );
    X_OPAD \RGB<5>/PAD (
      .PAD (RGB[5])
    );
    X_INV \RGB<5>/SRMUX (
      .I (N_RST),
      .O (\RGB[5]/SRNOT )
    );
    X_BUF \RGB<5>/OMUX (
      .I (rgb_int[5]),
      .O (\RGB[5]/OD )
    );
    X_BUF \C_RGB<5> (
      .I (N_RGB[5]),
      .O (\RGB[5]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<5>_218 (
      .I (\RGB[5]/OUTBUF_GTS_TRI ),
      .O (RGB[5]),
      .CTL (\C_RGB[5]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<5> (
      .I (\RGB[5]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[5]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[5])
    );
    X_OR2 \RGB<5>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[5]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[5]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<10>/KEEPER (
      .O (\RGB[10]/KEEPER )
    );
    X_OPAD \RGB<10>/PAD (
      .PAD (RGB[10])
    );
    X_INV \RGB<10>/SRMUX (
      .I (N_RST),
      .O (\RGB[10]/SRNOT )
    );
    X_BUF \RGB<10>/OMUX (
      .I (rgb_int[10]),
      .O (\RGB[10]/OD )
    );
    X_BUF \C_RGB<10> (
      .I (N_RGB[10]),
      .O (\RGB[10]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<10>_219 (
      .I (\RGB[10]/OUTBUF_GTS_TRI ),
      .O (RGB[10]),
      .CTL (\C_RGB[10]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<10> (
      .I (\RGB[10]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[10]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[10])
    );
    X_OR2 \RGB<10>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[10]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[10]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<6>/KEEPER (
      .O (\RGB[6]/KEEPER )
    );
    X_OPAD \RGB<6>/PAD (
      .PAD (RGB[6])
    );
    X_INV \RGB<6>/SRMUX (
      .I (N_RST),
      .O (\RGB[6]/SRNOT )
    );
    X_BUF \C_RGB<6> (
      .I (N_RGB[6]),
      .O (\RGB[6]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<6>_220 (
      .I (\RGB[6]/OUTBUF_GTS_TRI ),
      .O (RGB[6]),
      .CTL (\C_RGB[6]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<6> (
      .I (rgb_int[6]),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[6]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[6])
    );
    X_OR2 \RGB<6>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[6]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[6]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<11>/KEEPER (
      .O (\RGB[11]/KEEPER )
    );
    X_OPAD \RGB<11>/PAD (
      .PAD (RGB[11])
    );
    X_INV \RGB<11>/SRMUX (
      .I (N_RST),
      .O (\RGB[11]/SRNOT )
    );
    X_BUF \RGB<11>/OMUX (
      .I (rgb_int[11]),
      .O (\RGB[11]/OD )
    );
    X_BUF \C_RGB<11> (
      .I (N_RGB[11]),
      .O (\RGB[11]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<11>_221 (
      .I (\RGB[11]/OUTBUF_GTS_TRI ),
      .O (RGB[11]),
      .CTL (\C_RGB[11]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<11> (
      .I (\RGB[11]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[11]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[11])
    );
    X_OR2 \RGB<11>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[11]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[11]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<12>/KEEPER (
      .O (\RGB[12]/KEEPER )
    );
    X_OPAD \RGB<12>/PAD (
      .PAD (RGB[12])
    );
    X_INV \RGB<12>/SRMUX (
      .I (N_RST),
      .O (\RGB[12]/SRNOT )
    );
    X_BUF \RGB<12>/OMUX (
      .I (rgb_int[12]),
      .O (\RGB[12]/OD )
    );
    X_BUF \C_RGB<12> (
      .I (N_RGB[12]),
      .O (\RGB[12]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<12>_222 (
      .I (\RGB[12]/OUTBUF_GTS_TRI ),
      .O (RGB[12]),
      .CTL (\C_RGB[12]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<12> (
      .I (\RGB[12]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[12]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[12])
    );
    X_OR2 \RGB<12>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[12]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[12]/OFF/ASYNC_FF_GSR_OR )
    );
    X_KEEPER \RGB<13>/KEEPER (
      .O (\RGB[13]/KEEPER )
    );
    X_OPAD \RGB<13>/PAD (
      .PAD (RGB[13])
    );
    X_INV \RGB<13>/SRMUX (
      .I (N_RST),
      .O (\RGB[13]/SRNOT )
    );
    X_BUF \RGB<13>/OMUX (
      .I (rgb_int[13]),
      .O (\RGB[13]/OD )
    );
    X_BUF \C_RGB<13> (
      .I (N_RGB[13]),
      .O (\RGB[13]/OUTBUF_GTS_TRI )
    );
    X_TRI \C_RGB<13>_223 (
      .I (\RGB[13]/OUTBUF_GTS_TRI ),
      .O (RGB[13]),
      .CTL (\C_RGB[13]_2_INV )
    );
    X_FF \crt_out_reg/rgb_out_reg<13> (
      .I (\RGB[13]/OD ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\RGB[13]/OFF/ASYNC_FF_GSR_OR ),
      .O (N_RGB[13])
    );
    X_OR2 \RGB<13>/OFF/ASYNC_FF_GSR_OR (
      .I0 (\RGB[13]/SRNOT ),
      .I1 (GSR),
      .O (\RGB[13]/OFF/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[25]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<24> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [24]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [24])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<25> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [25]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [25])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[17]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<16> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [16]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [16])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<17> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [17]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [17])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<25>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[25]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<24> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [24]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [24])
    );
    X_OR2 \CRT/pix_start_addr<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[25]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<25> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [25]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [25])
    );
    X_OR2 \CRT/pix_start_addr<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[25]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[25]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \CRT/pix_start_addr<17>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[17]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<16> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [16]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [16])
    );
    X_OR2 \CRT/pix_start_addr<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[17]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<17> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [17]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [17])
    );
    X_OR2 \CRT/pix_start_addr<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[17]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[17]/FFX/ASYNC_FF_GSR_OR )
    );
    X_INV \bridge/pci_target_unit/pcit_if_bc_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_bc_out[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_bc_reg<2> (
      .I (\bridge/in_reg_cbe_out [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_bc_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_bc_out [2])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_bc_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_bc_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_bc_reg<3> (
      .I (\bridge/in_reg_cbe_out [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_bc_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_bc_out [3])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_bc_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_bc_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_bc_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_target_unit/pci_target_if/C5316/C2/C1/C0 .INIT = 16'hBB88;
    X_LUT4 \bridge/pci_target_unit/pci_target_if/C5316/C2/C1/C0 (
      .ADR0 (\bridge/pci_target_unit/pci_target_if/n_1335 ),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/conf_addr_out [0]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/n_1352 ),
      .O (\bridge/pci_target_unit/pci_target_if/C5316/C2/N8 )
    );
    defparam \bridge/pci_target_unit/pci_target_if/C5316/C2/C0/C0 .INIT = 16'hF0CC;
    X_LUT4 \bridge/pci_target_unit/pci_target_if/C5316/C2/C0/C0 (
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/pci_target_if/n_1317 ),
      .ADR2 (\bridge/pci_target_unit/pci_target_if/n_1298 ),
      .ADR3 (\bridge/pci_target_unit/pci_target_if/conf_addr_out [0]),
      .O (\bridge/pci_target_unit/pci_target_if/C5316/C2/N7 )
    );
    X_MUX2 \bridge/pci_target_unit/pci_target_if/C5316/C2/C2 (
      .IA (\bridge/pci_target_unit/pci_target_if/C5316/C2/N8 ),
      .IB (\bridge/pci_target_unit/pci_target_if/C5316/C2/N7 ),
      .SEL (\bridge/pci_target_unit/pci_target_if/conf_addr_out [1]),
      .O (\bridge/pci_target_unit/pci_target_if/N5157/F5MUX )
    );
    X_BUF \bridge/pci_target_unit/pci_target_if/N5157/XUSED (
      .I (\bridge/pci_target_unit/pci_target_if/N5157/F5MUX ),
      .O (\bridge/pci_target_unit/pci_target_if/N5157 )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C4/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C3/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C4/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C3/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3384/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3384/G (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3384/F .INIT = 16'hCCCC;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3384/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C3/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ONE ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C3/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ONE ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C3/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ZERO_224 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3384/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3385 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3384/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3384 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3384/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C4/C1/O )
    );
    X_ONE \bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ONE_225 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3384/LOGIC_ONE )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C6/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C5/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C6/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C5/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3386/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3386/G (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3386/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3386/F (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C5/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C4/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C5/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C4/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C5/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3386/LOGIC_ZERO_226 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3386/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3387 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3386/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3386 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3386/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3386/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C6/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C8/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C7/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C8/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C7/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3388/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3388/G (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3388/F .INIT = 16'hCCCC;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3388/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [6]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C7/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C6/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C7/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C6/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C7/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3388/LOGIC_ZERO_227 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3388/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3389 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3388/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3388 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3388/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3388/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C8/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C10/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C9/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C10/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C9/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3390/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3390/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [9]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3390/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3390/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [8]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C9/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C8/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C9/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C8/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C9/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3390/LOGIC_ZERO_228 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3390/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3391 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3390/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3390 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3390/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3390/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C10/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C12/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C11/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C12/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C11/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3392/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3392/G (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [11]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3392/F .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3392/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [10]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C11/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C10/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C11/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C10/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C11/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3392/LOGIC_ZERO_229 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3392/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3393 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3392/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3392 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3392/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3392/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C12/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C14/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C13/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C14/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C13/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3394/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3394/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [13]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3394/F .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3394/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [12]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C13/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C12/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C13/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C12/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C13/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3394/LOGIC_ZERO_230 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3394/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3395 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3394/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3394 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3394/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3394/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C14/C1/O )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[27]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<26> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [26]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [26])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<27> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [27]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [27])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C16/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C15/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C16/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C15/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3396/G .INIT = 16'hCCCC;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3396/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [15]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3396/F .INIT = 16'hCCCC;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3396/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [14]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C15/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C14/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C15/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C14/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C15/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3396/LOGIC_ZERO_231 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3396/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3397 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3396/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3396 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3396/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3396/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C16/C1/O )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[19]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<18> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [18]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [18])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<19> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [19]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [19])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C18/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C17/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C18/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C17/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3398/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3398/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [17]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3398/F .INIT = 16'hCCCC;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3398/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [16]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C17/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C16/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C17/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C16/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C17/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3398/LOGIC_ZERO_232 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3398/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3399 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3398/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3398 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3398/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3398/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C18/C1/O )
    );
    defparam \CRT/pix_start_addr<27>/F .INIT = 16'h0000;
    X_LUT4 \CRT/pix_start_addr<27>/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/pix_start_addr[27]/FROM )
    );
    X_INV \CRT/pix_start_addr<27>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[27]/SRNOT )
    );
    X_BUF \CRT/pix_start_addr<27>/XUSED (
      .I (\CRT/pix_start_addr[27]/FROM ),
      .O (GLOBAL_LOGIC0_1)
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<26> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [26]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [26])
    );
    X_OR2 \CRT/pix_start_addr<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[27]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<27> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [27]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [27])
    );
    X_OR2 \CRT/pix_start_addr<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[27]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[27]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C20/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C19/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C20/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C19/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3400/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3400/G (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [19]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3400/F .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3400/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [18]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C19/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C18/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C19/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C18/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C19/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3400/LOGIC_ZERO_233 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3400/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3401 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3400/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3400 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3400/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3400/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C20/C1/O )
    );
    X_INV \CRT/pix_start_addr<19>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[19]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<18> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [18]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [18])
    );
    X_OR2 \CRT/pix_start_addr<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[19]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<19> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [19]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [19])
    );
    X_OR2 \CRT/pix_start_addr<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[19]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[19]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C22/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C21/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C22/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C21/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3402/G .INIT = 16'hCCCC;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3402/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/pcim_if_address_out [21]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3402/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3402/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [20]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C21/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C20/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C21/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C20/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C21/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3402/LOGIC_ZERO_234 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3402/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3403 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3402/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3402 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3402/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3402/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C22/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C24/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C23/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C24/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C23/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3404/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3404/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [23]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3404/F .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3404/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [22]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C23/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C22/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C23/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C22/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C23/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3404/LOGIC_ZERO_235 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3404/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3405 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3404/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3404 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3404/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3404/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C24/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C26/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C25/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C26/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C25/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3406/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3406/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [25]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3406/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3406/F (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [24]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C25/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C24/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C25/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C24/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C25/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3406/LOGIC_ZERO_236 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3406/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3407 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3406/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3406 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3406/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3406/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C26/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C28/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C27/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C28/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C27/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3408/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3408/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [27]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3408/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3408/F (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [26]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C27/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C26/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C27/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C26/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C27/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3408/LOGIC_ZERO_237 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3408/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3409 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3408/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3408 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3408/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3408/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C28/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C30/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C29/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C30/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C29/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/GROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3410/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3410/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [29]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/GROM )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3410/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3410/F (
      .ADR0 (\bridge/wishbone_slave_unit/pcim_if_address_out [28]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C29/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C28/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C29/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C28/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C29/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3410/LOGIC_ZERO_238 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3410/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3411 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3410/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3410 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3410/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3410/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C30/C1/O )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[29]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<28> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [28]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [28])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<29> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [29]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [29])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C32/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C31/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pcim_if_address_out[31]_rt ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/XORG )
    );
    defparam \bridge/wishbone_slave_unit/pcim_if_address_out<31>_rt .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/pcim_if_address_out<31>_rt (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pcim_if_address_out [31]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pcim_if_address_out[31]_rt )
    );
    defparam \bridge/wishbone_slave_unit/pci_initiator_if/N3412/F .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/pci_initiator_if/N3412/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/pcim_if_address_out [30]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C31/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C30/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3274/C31/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C30/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/FROM ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3274/C31/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3412/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3413 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3412/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3412 )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3412/LOGIC_ZERO_239 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3412/LOGIC_ZERO )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C4/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C3/C1/O ),
      .I1 (\CRT/ssvga_fifo/N738/GROM ),
      .O (\CRT/ssvga_fifo/N738/XORG )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C4/C1 (
      .IA (\CRT/ssvga_fifo/N738/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C748/C3/C1/O ),
      .SEL (\CRT/ssvga_fifo/N738/GROM ),
      .O (\CRT/ssvga_fifo/N738/CYMUXG )
    );
    defparam \CRT/ssvga_fifo/N738/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_fifo/N738/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr_plus1 [1]),
      .O (\CRT/ssvga_fifo/N738/GROM )
    );
    defparam \CRT/ssvga_fifo/N738/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/N738/F (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [0]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N738/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C3/C0 (
      .I0 (\CRT/ssvga_fifo/N738/LOGIC_ONE ),
      .I1 (\CRT/ssvga_fifo/N738/FROM ),
      .O (\CRT/ssvga_fifo/N738/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C3/C1 (
      .IA (\CRT/ssvga_fifo/N738/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/N738/LOGIC_ONE ),
      .SEL (\CRT/ssvga_fifo/N738/FROM ),
      .O (\CRT/ssvga_fifo/C748/C3/C1/O )
    );
    X_ZERO \CRT/ssvga_fifo/N738/LOGIC_ZERO_240 (
      .O (\CRT/ssvga_fifo/N738/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_fifo/N738/YUSED (
      .I (\CRT/ssvga_fifo/N738/XORG ),
      .O (\CRT/ssvga_fifo/N739 )
    );
    X_BUF \CRT/ssvga_fifo/N738/XUSED (
      .I (\CRT/ssvga_fifo/N738/XORF ),
      .O (\CRT/ssvga_fifo/N738 )
    );
    X_BUF \CRT/ssvga_fifo/N738/COUTUSED (
      .I (\CRT/ssvga_fifo/N738/CYMUXG ),
      .O (\CRT/ssvga_fifo/C748/C4/C1/O )
    );
    X_ONE \CRT/ssvga_fifo/N738/LOGIC_ONE_241 (
      .O (\CRT/ssvga_fifo/N738/LOGIC_ONE )
    );
    X_INV \CRT/pix_start_addr<29>/SRMUX (
      .I (N_RST),
      .O (\CRT/pix_start_addr[29]/SRNOT )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<28> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [28]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [28])
    );
    X_OR2 \CRT/pix_start_addr<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[29]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \CRT/ssvga_wbs_if/pix_start_addr_reg<29> (
      .I (\bridge/pci_target_unit/fifos_pciw_addr_data_out [29]),
      .CLK (CLK_BUFGPed),
      .CE (N12120),
      .SET (GND),
      .RST (\CRT/pix_start_addr[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\CRT/pix_start_addr [29])
    );
    X_OR2 \CRT/pix_start_addr<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\CRT/pix_start_addr[29]/SRNOT ),
      .I1 (GSR),
      .O (\CRT/pix_start_addr[29]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C6/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C5/C1/O ),
      .I1 (\CRT/ssvga_fifo/N740/GROM ),
      .O (\CRT/ssvga_fifo/N740/XORG )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C6/C1 (
      .IA (\CRT/ssvga_fifo/N740/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C748/C5/C1/O ),
      .SEL (\CRT/ssvga_fifo/N740/GROM ),
      .O (\CRT/ssvga_fifo/N740/CYMUXG )
    );
    defparam \CRT/ssvga_fifo/N740/G .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_fifo/N740/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr_plus1 [3]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N740/GROM )
    );
    defparam \CRT/ssvga_fifo/N740/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_fifo/N740/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/rd_ptr_plus1 [2]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N740/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C5/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C4/C1/O ),
      .I1 (\CRT/ssvga_fifo/N740/FROM ),
      .O (\CRT/ssvga_fifo/N740/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C5/C1 (
      .IA (\CRT/ssvga_fifo/N740/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C748/C4/C1/O ),
      .SEL (\CRT/ssvga_fifo/N740/FROM ),
      .O (\CRT/ssvga_fifo/C748/C5/C1/O )
    );
    X_ZERO \CRT/ssvga_fifo/N740/LOGIC_ZERO_242 (
      .O (\CRT/ssvga_fifo/N740/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_fifo/N740/YUSED (
      .I (\CRT/ssvga_fifo/N740/XORG ),
      .O (\CRT/ssvga_fifo/N741 )
    );
    X_BUF \CRT/ssvga_fifo/N740/XUSED (
      .I (\CRT/ssvga_fifo/N740/XORF ),
      .O (\CRT/ssvga_fifo/N740 )
    );
    X_BUF \CRT/ssvga_fifo/N740/COUTUSED (
      .I (\CRT/ssvga_fifo/N740/CYMUXG ),
      .O (\CRT/ssvga_fifo/C748/C6/C1/O )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C8/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C7/C1/O ),
      .I1 (\CRT/ssvga_fifo/N742/GROM ),
      .O (\CRT/ssvga_fifo/N742/XORG )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C8/C1 (
      .IA (\CRT/ssvga_fifo/N742/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C748/C7/C1/O ),
      .SEL (\CRT/ssvga_fifo/N742/GROM ),
      .O (\CRT/ssvga_fifo/N742/CYMUXG )
    );
    defparam \CRT/ssvga_fifo/N742/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_fifo/N742/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr_plus1 [5]),
      .O (\CRT/ssvga_fifo/N742/GROM )
    );
    defparam \CRT/ssvga_fifo/N742/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/N742/F (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [4]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N742/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C7/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C6/C1/O ),
      .I1 (\CRT/ssvga_fifo/N742/FROM ),
      .O (\CRT/ssvga_fifo/N742/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C7/C1 (
      .IA (\CRT/ssvga_fifo/N742/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C748/C6/C1/O ),
      .SEL (\CRT/ssvga_fifo/N742/FROM ),
      .O (\CRT/ssvga_fifo/C748/C7/C1/O )
    );
    X_ZERO \CRT/ssvga_fifo/N742/LOGIC_ZERO_243 (
      .O (\CRT/ssvga_fifo/N742/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_fifo/N742/YUSED (
      .I (\CRT/ssvga_fifo/N742/XORG ),
      .O (\CRT/ssvga_fifo/N743 )
    );
    X_BUF \CRT/ssvga_fifo/N742/XUSED (
      .I (\CRT/ssvga_fifo/N742/XORF ),
      .O (\CRT/ssvga_fifo/N742 )
    );
    X_BUF \CRT/ssvga_fifo/N742/COUTUSED (
      .I (\CRT/ssvga_fifo/N742/CYMUXG ),
      .O (\CRT/ssvga_fifo/C748/C8/C1/O )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C10/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C9/C1/O ),
      .I1 (\CRT/ssvga_fifo/N744/GROM ),
      .O (\CRT/ssvga_fifo/N744/XORG )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C10/C1 (
      .IA (\CRT/ssvga_fifo/N744/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C748/C9/C1/O ),
      .SEL (\CRT/ssvga_fifo/N744/GROM ),
      .O (\CRT/ssvga_fifo/N744/CYMUXG )
    );
    defparam \CRT/ssvga_fifo/N744/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/N744/G (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [7]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N744/GROM )
    );
    defparam \CRT/ssvga_fifo/N744/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/N744/F (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [6]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N744/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C9/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C8/C1/O ),
      .I1 (\CRT/ssvga_fifo/N744/FROM ),
      .O (\CRT/ssvga_fifo/N744/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C9/C1 (
      .IA (\CRT/ssvga_fifo/N744/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C748/C8/C1/O ),
      .SEL (\CRT/ssvga_fifo/N744/FROM ),
      .O (\CRT/ssvga_fifo/C748/C9/C1/O )
    );
    X_ZERO \CRT/ssvga_fifo/N744/LOGIC_ZERO_244 (
      .O (\CRT/ssvga_fifo/N744/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_fifo/N744/YUSED (
      .I (\CRT/ssvga_fifo/N744/XORG ),
      .O (\CRT/ssvga_fifo/N745 )
    );
    X_BUF \CRT/ssvga_fifo/N744/XUSED (
      .I (\CRT/ssvga_fifo/N744/XORF ),
      .O (\CRT/ssvga_fifo/N744 )
    );
    X_BUF \CRT/ssvga_fifo/N744/COUTUSED (
      .I (\CRT/ssvga_fifo/N744/CYMUXG ),
      .O (\CRT/ssvga_fifo/C748/C10/C1/O )
    );
    X_ONE \bridge/configuration/pci_error_rty_exp_set/LOGIC_ONE_245 (
      .O (\bridge/configuration/pci_error_rty_exp_set/LOGIC_ONE )
    );
    X_FF \bridge/configuration/pci_err_cs_bit10_reg (
      .I (\bridge/configuration/pci_error_rty_exp_set/LOGIC_ONE ),
      .CLK (CLK_BUFGPed),
      .CE (N12312),
      .SET (GND),
      .RST (\bridge/configuration/pci_error_rty_exp_set/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/configuration/pci_error_rty_exp_set )
    );
    X_OR2 \bridge/configuration/pci_error_rty_exp_set/FFY/ASYNC_FF_GSR_OR_246 (
      .I0 (\bridge/configuration/delete_pci_err_cs_bit10 ),
      .I1 (GSR),
      .O (\bridge/configuration/pci_error_rty_exp_set/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C12/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C11/C1/O ),
      .I1 (\CRT/ssvga_fifo/rd_ptr_plus1[9]_rt ),
      .O (\CRT/ssvga_fifo/N746/XORG )
    );
    defparam \CRT/ssvga_fifo/rd_ptr_plus1<9>_rt .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/rd_ptr_plus1<9>_rt (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/rd_ptr_plus1 [9]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/rd_ptr_plus1[9]_rt )
    );
    defparam \CRT/ssvga_fifo/N746/F .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_fifo/N746/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_fifo/rd_ptr_plus1 [8]),
      .O (\CRT/ssvga_fifo/N746/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C748/C11/C0 (
      .I0 (\CRT/ssvga_fifo/C748/C10/C1/O ),
      .I1 (\CRT/ssvga_fifo/N746/FROM ),
      .O (\CRT/ssvga_fifo/N746/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C748/C11/C1 (
      .IA (\CRT/ssvga_fifo/N746/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C748/C10/C1/O ),
      .SEL (\CRT/ssvga_fifo/N746/FROM ),
      .O (\CRT/ssvga_fifo/C748/C11/C1/O )
    );
    X_BUF \CRT/ssvga_fifo/N746/YUSED (
      .I (\CRT/ssvga_fifo/N746/XORG ),
      .O (\CRT/ssvga_fifo/N747 )
    );
    X_BUF \CRT/ssvga_fifo/N746/XUSED (
      .I (\CRT/ssvga_fifo/N746/XORF ),
      .O (\CRT/ssvga_fifo/N746 )
    );
    X_ZERO \CRT/ssvga_fifo/N746/LOGIC_ZERO_247 (
      .O (\CRT/ssvga_fifo/N746/LOGIC_ZERO )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C4/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C3/C1/O ),
      .I1 (N12625),
      .O (\CRT/ssvga_wbm_if/N1515/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C4/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [1]),
      .IB (\CRT/ssvga_wbm_if/C1472/C3/C1/O ),
      .SEL (N12625),
      .O (\CRT/ssvga_wbm_if/N1515/CYMUXG )
    );
    defparam C19125.INIT = 16'h5555;
    X_LUT4 C19125(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [1]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12625)
    );
    defparam C19126.INIT = 16'h5555;
    X_LUT4 C19126(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [0]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12642)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C3/C0 (
      .I0 (\CRT/ssvga_wbm_if/N1515/LOGIC_ZERO ),
      .I1 (N12642),
      .O (\CRT/ssvga_wbm_if/N1515/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C3/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [0]),
      .IB (\CRT/ssvga_wbm_if/N1515/LOGIC_ZERO ),
      .SEL (N12642),
      .O (\CRT/ssvga_wbm_if/C1472/C3/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1515/YUSED (
      .I (\CRT/ssvga_wbm_if/N1515/XORG ),
      .O (\CRT/ssvga_wbm_if/N1516 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1515/XUSED (
      .I (\CRT/ssvga_wbm_if/N1515/XORF ),
      .O (\CRT/ssvga_wbm_if/N1515 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1515/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1515/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1472/C4/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1515/LOGIC_ZERO_248 (
      .O (\CRT/ssvga_wbm_if/N1515/LOGIC_ZERO )
    );
    X_INV \bridge/pci_target_unit/pci_target_if/bckp_trdy_reg/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pci_target_if/bckp_trdy_reg/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/bckp_trdy_reg_reg (
      .I (\bridge/out_bckp_trdy_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/pci_target_if/bckp_trdy_reg/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pci_target_if/bckp_trdy_reg )
    );
    X_OR2
     \bridge/pci_target_unit/pci_target_if/bckp_trdy_reg/FFY/ASYNC_FF_GSR_OR_249 (
      .I0 (\bridge/pci_target_unit/pci_target_if/bckp_trdy_reg/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/pci_target_if/bckp_trdy_reg/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C6/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C5/C1/O ),
      .I1 (N12619),
      .O (\CRT/ssvga_wbm_if/N1517/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C6/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [3]),
      .IB (\CRT/ssvga_wbm_if/C1472/C5/C1/O ),
      .SEL (N12619),
      .O (\CRT/ssvga_wbm_if/N1517/CYMUXG )
    );
    defparam C19123.INIT = 16'h5555;
    X_LUT4 C19123(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12619)
    );
    defparam C19124.INIT = 16'h5555;
    X_LUT4 C19124(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [2]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12650)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C5/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C4/C1/O ),
      .I1 (N12650),
      .O (\CRT/ssvga_wbm_if/N1517/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C5/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [2]),
      .IB (\CRT/ssvga_wbm_if/C1472/C4/C1/O ),
      .SEL (N12650),
      .O (\CRT/ssvga_wbm_if/C1472/C5/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1517/YUSED (
      .I (\CRT/ssvga_wbm_if/N1517/XORG ),
      .O (\CRT/ssvga_wbm_if/N1518 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1517/XUSED (
      .I (\CRT/ssvga_wbm_if/N1517/XORF ),
      .O (\CRT/ssvga_wbm_if/N1517 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1517/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1517/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1472/C6/C1/O )
    );
    X_INV \bridge/conf_cache_line_size_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_cache_line_size_out[1]/SRNOT )
    );
    X_FF \bridge/configuration/cache_line_size_reg_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C284/N39 ),
      .SET (GND),
      .RST (\bridge/conf_cache_line_size_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_cache_line_size_out [0])
    );
    X_OR2 \bridge/conf_cache_line_size_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_cache_line_size_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_cache_line_size_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cache_line_size_reg_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C284/N39 ),
      .SET (GND),
      .RST (\bridge/conf_cache_line_size_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_cache_line_size_out [1])
    );
    X_OR2 \bridge/conf_cache_line_size_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_cache_line_size_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_cache_line_size_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C8/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C7/C1/O ),
      .I1 (N12623),
      .O (\CRT/ssvga_wbm_if/N1519/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C8/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [5]),
      .IB (\CRT/ssvga_wbm_if/C1472/C7/C1/O ),
      .SEL (N12623),
      .O (\CRT/ssvga_wbm_if/N1519/CYMUXG )
    );
    defparam C19121.INIT = 16'h5555;
    X_LUT4 C19121(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12623)
    );
    defparam C19122.INIT = 16'h5555;
    X_LUT4 C19122(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12646)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C7/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C6/C1/O ),
      .I1 (N12646),
      .O (\CRT/ssvga_wbm_if/N1519/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C7/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [4]),
      .IB (\CRT/ssvga_wbm_if/C1472/C6/C1/O ),
      .SEL (N12646),
      .O (\CRT/ssvga_wbm_if/C1472/C7/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1519/YUSED (
      .I (\CRT/ssvga_wbm_if/N1519/XORG ),
      .O (\CRT/ssvga_wbm_if/N1520 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1519/XUSED (
      .I (\CRT/ssvga_wbm_if/N1519/XORF ),
      .O (\CRT/ssvga_wbm_if/N1519 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1519/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1519/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1472/C8/C1/O )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C10/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C9/C1/O ),
      .I1 (N12621),
      .O (\CRT/ssvga_wbm_if/N1521/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C10/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [7]),
      .IB (\CRT/ssvga_wbm_if/C1472/C9/C1/O ),
      .SEL (N12621),
      .O (\CRT/ssvga_wbm_if/N1521/CYMUXG )
    );
    defparam C19119.INIT = 16'h5555;
    X_LUT4 C19119(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12621)
    );
    defparam C19120.INIT = 16'h5555;
    X_LUT4 C19120(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [6]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12648)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C9/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C8/C1/O ),
      .I1 (N12648),
      .O (\CRT/ssvga_wbm_if/N1521/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C9/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [6]),
      .IB (\CRT/ssvga_wbm_if/C1472/C8/C1/O ),
      .SEL (N12648),
      .O (\CRT/ssvga_wbm_if/C1472/C9/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1521/YUSED (
      .I (\CRT/ssvga_wbm_if/N1521/XORG ),
      .O (\CRT/ssvga_wbm_if/N1522 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1521/XUSED (
      .I (\CRT/ssvga_wbm_if/N1521/XORF ),
      .O (\CRT/ssvga_wbm_if/N1521 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1521/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1521/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1472/C10/C1/O )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C12/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C11/C1/O ),
      .I1 (N12644),
      .O (\CRT/ssvga_wbm_if/N1523/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C12/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [9]),
      .IB (\CRT/ssvga_wbm_if/C1472/C11/C1/O ),
      .SEL (N12644),
      .O (\CRT/ssvga_wbm_if/N1523/CYMUXG )
    );
    defparam C19117.INIT = 16'h5555;
    X_LUT4 C19117(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [9]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12644)
    );
    defparam C19118.INIT = 16'h5555;
    X_LUT4 C19118(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [8]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12627)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C11/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C10/C1/O ),
      .I1 (N12627),
      .O (\CRT/ssvga_wbm_if/N1523/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C11/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [8]),
      .IB (\CRT/ssvga_wbm_if/C1472/C10/C1/O ),
      .SEL (N12627),
      .O (\CRT/ssvga_wbm_if/C1472/C11/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1523/YUSED (
      .I (\CRT/ssvga_wbm_if/N1523/XORG ),
      .O (\CRT/ssvga_wbm_if/N1524 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1523/XUSED (
      .I (\CRT/ssvga_wbm_if/N1523/XORF ),
      .O (\CRT/ssvga_wbm_if/N1523 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1523/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1523/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1472/C12/C1/O )
    );
    X_INV \bridge/conf_cache_line_size_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_cache_line_size_out[3]/SRNOT )
    );
    X_FF \bridge/configuration/cache_line_size_reg_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C284/N39 ),
      .SET (GND),
      .RST (\bridge/conf_cache_line_size_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_cache_line_size_out [2])
    );
    X_OR2 \bridge/conf_cache_line_size_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_cache_line_size_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_cache_line_size_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cache_line_size_reg_reg<3> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C284/N39 ),
      .SET (GND),
      .RST (\bridge/conf_cache_line_size_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_cache_line_size_out [3])
    );
    X_OR2 \bridge/conf_cache_line_size_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_cache_line_size_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_cache_line_size_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C14/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C13/C1/O ),
      .I1 (N12631),
      .O (\CRT/ssvga_wbm_if/N1525/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C14/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [11]),
      .IB (\CRT/ssvga_wbm_if/C1472/C13/C1/O ),
      .SEL (N12631),
      .O (\CRT/ssvga_wbm_if/N1525/CYMUXG )
    );
    defparam C19115.INIT = 16'h5555;
    X_LUT4 C19115(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [11]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12631)
    );
    defparam C19116.INIT = 16'h5555;
    X_LUT4 C19116(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [10]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12638)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C13/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C12/C1/O ),
      .I1 (N12638),
      .O (\CRT/ssvga_wbm_if/N1525/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C13/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [10]),
      .IB (\CRT/ssvga_wbm_if/C1472/C12/C1/O ),
      .SEL (N12638),
      .O (\CRT/ssvga_wbm_if/C1472/C13/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1525/YUSED (
      .I (\CRT/ssvga_wbm_if/N1525/XORG ),
      .O (\CRT/ssvga_wbm_if/N1526 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1525/XUSED (
      .I (\CRT/ssvga_wbm_if/N1525/XORF ),
      .O (\CRT/ssvga_wbm_if/N1525 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1525/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1525/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1472/C14/C1/O )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C16/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C15/C1/O ),
      .I1 (N12633),
      .O (\CRT/ssvga_wbm_if/N1527/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C16/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [13]),
      .IB (\CRT/ssvga_wbm_if/C1472/C15/C1/O ),
      .SEL (N12633),
      .O (\CRT/ssvga_wbm_if/N1527/CYMUXG )
    );
    defparam C19113.INIT = 16'h5555;
    X_LUT4 C19113(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [13]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12633)
    );
    defparam C19114.INIT = 16'h5555;
    X_LUT4 C19114(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [12]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12636)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C15/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C14/C1/O ),
      .I1 (N12636),
      .O (\CRT/ssvga_wbm_if/N1527/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C15/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [12]),
      .IB (\CRT/ssvga_wbm_if/C1472/C14/C1/O ),
      .SEL (N12636),
      .O (\CRT/ssvga_wbm_if/C1472/C15/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1527/YUSED (
      .I (\CRT/ssvga_wbm_if/N1527/XORG ),
      .O (\CRT/ssvga_wbm_if/N1528 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1527/XUSED (
      .I (\CRT/ssvga_wbm_if/N1527/XORF ),
      .O (\CRT/ssvga_wbm_if/N1527 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1527/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1527/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1472/C16/C1/O )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C18/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C17/C1/O ),
      .I1 (N12629),
      .O (\CRT/ssvga_wbm_if/N1529/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C18/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [15]),
      .IB (\CRT/ssvga_wbm_if/C1472/C17/C1/O ),
      .SEL (N12629),
      .O (\CRT/ssvga_wbm_if/N1529/CYMUXG )
    );
    defparam C19111.INIT = 16'h5555;
    X_LUT4 C19111(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [15]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12629)
    );
    defparam C19112.INIT = 16'h5555;
    X_LUT4 C19112(
      .ADR0 (\CRT/ssvga_wbm_if/vmaddr_r [14]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12640)
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1472/C17/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1472/C16/C1/O ),
      .I1 (N12640),
      .O (\CRT/ssvga_wbm_if/N1529/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1472/C17/C1 (
      .IA (\CRT/ssvga_wbm_if/vmaddr_r [14]),
      .IB (\CRT/ssvga_wbm_if/C1472/C16/C1/O ),
      .SEL (N12640),
      .O (\CRT/ssvga_wbm_if/C1472/C17/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1529/YUSED (
      .I (\CRT/ssvga_wbm_if/N1529/XORG ),
      .O (\CRT/ssvga_wbm_if/N1530 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1529/XUSED (
      .I (\CRT/ssvga_wbm_if/N1529/XORF ),
      .O (\CRT/ssvga_wbm_if/N1529 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1529/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1529/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1472/C18/C1/O )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_XOR2 \CRT/ssvga_fifo/C749/C4/C0 (
      .I0 (\CRT/ssvga_fifo/C749/C3/C1/O ),
      .I1 (\CRT/ssvga_fifo/N800/GROM ),
      .O (\CRT/ssvga_fifo/N800/XORG )
    );
    X_MUX2 \CRT/ssvga_fifo/C749/C4/C1 (
      .IA (\CRT/ssvga_fifo/N800/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C749/C3/C1/O ),
      .SEL (\CRT/ssvga_fifo/N800/GROM ),
      .O (\CRT/ssvga_fifo/N800/CYMUXG )
    );
    defparam \CRT/ssvga_fifo/N800/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/N800/G (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [1]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N800/GROM )
    );
    defparam \CRT/ssvga_fifo/N800/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_fifo/N800/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [0]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N800/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C749/C3/C0 (
      .I0 (\CRT/ssvga_fifo/N800/LOGIC_ONE ),
      .I1 (\CRT/ssvga_fifo/N800/FROM ),
      .O (\CRT/ssvga_fifo/N800/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C749/C3/C1 (
      .IA (\CRT/ssvga_fifo/N800/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/N800/LOGIC_ONE ),
      .SEL (\CRT/ssvga_fifo/N800/FROM ),
      .O (\CRT/ssvga_fifo/C749/C3/C1/O )
    );
    X_ZERO \CRT/ssvga_fifo/N800/LOGIC_ZERO_250 (
      .O (\CRT/ssvga_fifo/N800/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_fifo/N800/YUSED (
      .I (\CRT/ssvga_fifo/N800/XORG ),
      .O (\CRT/ssvga_fifo/N801 )
    );
    X_BUF \CRT/ssvga_fifo/N800/XUSED (
      .I (\CRT/ssvga_fifo/N800/XORF ),
      .O (\CRT/ssvga_fifo/N800 )
    );
    X_BUF \CRT/ssvga_fifo/N800/COUTUSED (
      .I (\CRT/ssvga_fifo/N800/CYMUXG ),
      .O (\CRT/ssvga_fifo/C749/C4/C1/O )
    );
    X_ONE \CRT/ssvga_fifo/N800/LOGIC_ONE_251 (
      .O (\CRT/ssvga_fifo/N800/LOGIC_ONE )
    );
    X_INV \bridge/conf_cache_line_size_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_cache_line_size_out[5]/SRNOT )
    );
    X_FF \bridge/configuration/cache_line_size_reg_reg<4> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C284/N39 ),
      .SET (GND),
      .RST (\bridge/conf_cache_line_size_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_cache_line_size_out [4])
    );
    X_OR2 \bridge/conf_cache_line_size_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_cache_line_size_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_cache_line_size_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cache_line_size_reg_reg<5> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C284/N39 ),
      .SET (GND),
      .RST (\bridge/conf_cache_line_size_out[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_cache_line_size_out [5])
    );
    X_OR2 \bridge/conf_cache_line_size_out<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_cache_line_size_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_cache_line_size_out[5]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_fifo/C749/C6/C0 (
      .I0 (\CRT/ssvga_fifo/C749/C5/C1/O ),
      .I1 (\CRT/ssvga_fifo/N802/GROM ),
      .O (\CRT/ssvga_fifo/N802/XORG )
    );
    X_MUX2 \CRT/ssvga_fifo/C749/C6/C1 (
      .IA (\CRT/ssvga_fifo/N802/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C749/C5/C1/O ),
      .SEL (\CRT/ssvga_fifo/N802/GROM ),
      .O (\CRT/ssvga_fifo/N802/CYMUXG )
    );
    defparam \CRT/ssvga_fifo/N802/G .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_fifo/N802/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [3]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N802/GROM )
    );
    defparam \CRT/ssvga_fifo/N802/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/N802/F (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N802/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C749/C5/C0 (
      .I0 (\CRT/ssvga_fifo/C749/C4/C1/O ),
      .I1 (\CRT/ssvga_fifo/N802/FROM ),
      .O (\CRT/ssvga_fifo/N802/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C749/C5/C1 (
      .IA (\CRT/ssvga_fifo/N802/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C749/C4/C1/O ),
      .SEL (\CRT/ssvga_fifo/N802/FROM ),
      .O (\CRT/ssvga_fifo/C749/C5/C1/O )
    );
    X_ZERO \CRT/ssvga_fifo/N802/LOGIC_ZERO_252 (
      .O (\CRT/ssvga_fifo/N802/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_fifo/N802/YUSED (
      .I (\CRT/ssvga_fifo/N802/XORG ),
      .O (\CRT/ssvga_fifo/N803 )
    );
    X_BUF \CRT/ssvga_fifo/N802/XUSED (
      .I (\CRT/ssvga_fifo/N802/XORF ),
      .O (\CRT/ssvga_fifo/N802 )
    );
    X_BUF \CRT/ssvga_fifo/N802/COUTUSED (
      .I (\CRT/ssvga_fifo/N802/CYMUXG ),
      .O (\CRT/ssvga_fifo/C749/C6/C1/O )
    );
    X_XOR2 \CRT/ssvga_fifo/C749/C8/C0 (
      .I0 (\CRT/ssvga_fifo/C749/C7/C1/O ),
      .I1 (\CRT/ssvga_fifo/N804/GROM ),
      .O (\CRT/ssvga_fifo/N804/XORG )
    );
    X_MUX2 \CRT/ssvga_fifo/C749/C8/C1 (
      .IA (\CRT/ssvga_fifo/N804/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C749/C7/C1/O ),
      .SEL (\CRT/ssvga_fifo/N804/GROM ),
      .O (\CRT/ssvga_fifo/N804/CYMUXG )
    );
    defparam \CRT/ssvga_fifo/N804/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/N804/G (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [5]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N804/GROM )
    );
    defparam \CRT/ssvga_fifo/N804/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_fifo/N804/F (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_fifo/wr_ptr_plus1 [4]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N804/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C749/C7/C0 (
      .I0 (\CRT/ssvga_fifo/C749/C6/C1/O ),
      .I1 (\CRT/ssvga_fifo/N804/FROM ),
      .O (\CRT/ssvga_fifo/N804/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C749/C7/C1 (
      .IA (\CRT/ssvga_fifo/N804/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C749/C6/C1/O ),
      .SEL (\CRT/ssvga_fifo/N804/FROM ),
      .O (\CRT/ssvga_fifo/C749/C7/C1/O )
    );
    X_ZERO \CRT/ssvga_fifo/N804/LOGIC_ZERO_253 (
      .O (\CRT/ssvga_fifo/N804/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_fifo/N804/YUSED (
      .I (\CRT/ssvga_fifo/N804/XORG ),
      .O (\CRT/ssvga_fifo/N805 )
    );
    X_BUF \CRT/ssvga_fifo/N804/XUSED (
      .I (\CRT/ssvga_fifo/N804/XORF ),
      .O (\CRT/ssvga_fifo/N804 )
    );
    X_BUF \CRT/ssvga_fifo/N804/COUTUSED (
      .I (\CRT/ssvga_fifo/N804/CYMUXG ),
      .O (\CRT/ssvga_fifo/C749/C8/C1/O )
    );
    X_XOR2 \CRT/ssvga_fifo/C749/C10/C0 (
      .I0 (\CRT/ssvga_fifo/C749/C9/C1/O ),
      .I1 (\CRT/ssvga_fifo/wr_ptr_plus1[7]_rt ),
      .O (\CRT/ssvga_fifo/N806/XORG )
    );
    defparam \CRT/ssvga_fifo/wr_ptr_plus1<7>_rt .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_fifo/wr_ptr_plus1<7>_rt (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [7]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/wr_ptr_plus1[7]_rt )
    );
    defparam \CRT/ssvga_fifo/N806/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_fifo/N806/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_fifo/wr_ptr_plus1 [6]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_fifo/N806/FROM )
    );
    X_XOR2 \CRT/ssvga_fifo/C749/C9/C0 (
      .I0 (\CRT/ssvga_fifo/C749/C8/C1/O ),
      .I1 (\CRT/ssvga_fifo/N806/FROM ),
      .O (\CRT/ssvga_fifo/N806/XORF )
    );
    X_MUX2 \CRT/ssvga_fifo/C749/C9/C1 (
      .IA (\CRT/ssvga_fifo/N806/LOGIC_ZERO ),
      .IB (\CRT/ssvga_fifo/C749/C8/C1/O ),
      .SEL (\CRT/ssvga_fifo/N806/FROM ),
      .O (\CRT/ssvga_fifo/C749/C9/C1/O )
    );
    X_BUF \CRT/ssvga_fifo/N806/YUSED (
      .I (\CRT/ssvga_fifo/N806/XORG ),
      .O (\CRT/ssvga_fifo/N807 )
    );
    X_BUF \CRT/ssvga_fifo/N806/XUSED (
      .I (\CRT/ssvga_fifo/N806/XORF ),
      .O (\CRT/ssvga_fifo/N806 )
    );
    X_ZERO \CRT/ssvga_fifo/N806/LOGIC_ZERO_254 (
      .O (\CRT/ssvga_fifo/N806/LOGIC_ZERO )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[4]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[4]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C4/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C3/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1235/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1235/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C4/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1235/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C3/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1235/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1235/CYMUXG )
    );
    defparam \bridge/pci_target_unit/del_sync/N1235/G .INIT = 16'hCCCC;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1235/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/comp_cycle_count [1]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1235/GROM )
    );
    defparam \bridge/pci_target_unit/del_sync/N1235/F .INIT = 16'hFF00;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1235/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/comp_cycle_count [0]),
      .O (\bridge/pci_target_unit/del_sync/N1235/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C3/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/N1235/LOGIC_ONE ),
      .I1 (\bridge/pci_target_unit/del_sync/N1235/FROM ),
      .O (\bridge/pci_target_unit/del_sync/N1235/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C3/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1235/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/N1235/LOGIC_ONE ),
      .SEL (\bridge/pci_target_unit/del_sync/N1235/FROM ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C3/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/del_sync/N1235/LOGIC_ZERO_255 (
      .O (\bridge/pci_target_unit/del_sync/N1235/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1235/YUSED (
      .I (\bridge/pci_target_unit/del_sync/N1235/XORG ),
      .O (\bridge/pci_target_unit/del_sync/N1236 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1235/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1235/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1235 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1235/COUTUSED (
      .I (\bridge/pci_target_unit/del_sync/N1235/CYMUXG ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C4/C1/O )
    );
    X_ONE \bridge/pci_target_unit/del_sync/N1235/LOGIC_ONE_256 (
      .O (\bridge/pci_target_unit/del_sync/N1235/LOGIC_ONE )
    );
    X_INV \bridge/conf_cache_line_size_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_cache_line_size_out[7]/SRNOT )
    );
    X_FF \bridge/configuration/cache_line_size_reg_reg<6> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C284/N39 ),
      .SET (GND),
      .RST (\bridge/conf_cache_line_size_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_cache_line_size_out [6])
    );
    X_OR2 \bridge/conf_cache_line_size_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_cache_line_size_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_cache_line_size_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/configuration/cache_line_size_reg_reg<7> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C284/N39 ),
      .SET (GND),
      .RST (\bridge/conf_cache_line_size_out[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_cache_line_size_out [7])
    );
    X_OR2 \bridge/conf_cache_line_size_out<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/conf_cache_line_size_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_cache_line_size_out[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C6/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C5/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1237/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1237/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C6/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1237/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C5/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1237/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1237/CYMUXG )
    );
    defparam \bridge/pci_target_unit/del_sync/N1237/G .INIT = 16'hCCCC;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1237/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/comp_cycle_count [3]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1237/GROM )
    );
    defparam \bridge/pci_target_unit/del_sync/N1237/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1237/F (
      .ADR0 (\bridge/pci_target_unit/del_sync/comp_cycle_count [2]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1237/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C5/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C4/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1237/FROM ),
      .O (\bridge/pci_target_unit/del_sync/N1237/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C5/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1237/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C4/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1237/FROM ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C5/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/del_sync/N1237/LOGIC_ZERO_257 (
      .O (\bridge/pci_target_unit/del_sync/N1237/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1237/YUSED (
      .I (\bridge/pci_target_unit/del_sync/N1237/XORG ),
      .O (\bridge/pci_target_unit/del_sync/N1238 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1237/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1237/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1237 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1237/COUTUSED (
      .I (\bridge/pci_target_unit/del_sync/N1237/CYMUXG ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C6/C1/O )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C8/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C7/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1239/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1239/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C8/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1239/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C7/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1239/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1239/CYMUXG )
    );
    defparam \bridge/pci_target_unit/del_sync/N1239/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1239/G (
      .ADR0 (\bridge/pci_target_unit/del_sync/comp_cycle_count [5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1239/GROM )
    );
    defparam \bridge/pci_target_unit/del_sync/N1239/F .INIT = 16'hCCCC;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1239/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/comp_cycle_count [4]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1239/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C7/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C6/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1239/FROM ),
      .O (\bridge/pci_target_unit/del_sync/N1239/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C7/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1239/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C6/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1239/FROM ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C7/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/del_sync/N1239/LOGIC_ZERO_258 (
      .O (\bridge/pci_target_unit/del_sync/N1239/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1239/YUSED (
      .I (\bridge/pci_target_unit/del_sync/N1239/XORG ),
      .O (\bridge/pci_target_unit/del_sync/N1240 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1239/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1239/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1239 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1239/COUTUSED (
      .I (\bridge/pci_target_unit/del_sync/N1239/CYMUXG ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C8/C1/O )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<0> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [0])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<1> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [1])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[1]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[1]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C10/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C9/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1241/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1241/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C10/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1241/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C9/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1241/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1241/CYMUXG )
    );
    defparam \bridge/pci_target_unit/del_sync/N1241/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1241/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_cycle_count [7]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1241/GROM )
    );
    defparam \bridge/pci_target_unit/del_sync/N1241/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1241/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_cycle_count [6]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1241/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C9/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C8/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1241/FROM ),
      .O (\bridge/pci_target_unit/del_sync/N1241/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C9/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1241/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C8/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1241/FROM ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C9/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/del_sync/N1241/LOGIC_ZERO_259 (
      .O (\bridge/pci_target_unit/del_sync/N1241/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1241/YUSED (
      .I (\bridge/pci_target_unit/del_sync/N1241/XORG ),
      .O (\bridge/pci_target_unit/del_sync/N1242 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1241/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1241/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1241 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1241/COUTUSED (
      .I (\bridge/pci_target_unit/del_sync/N1241/CYMUXG ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C10/C1/O )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C12/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C11/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1243/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1243/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C12/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1243/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C11/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1243/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1243/CYMUXG )
    );
    defparam \bridge/pci_target_unit/del_sync/N1243/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1243/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_cycle_count [9]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1243/GROM )
    );
    defparam \bridge/pci_target_unit/del_sync/N1243/F .INIT = 16'hFF00;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1243/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/comp_cycle_count [8]),
      .O (\bridge/pci_target_unit/del_sync/N1243/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C11/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C10/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1243/FROM ),
      .O (\bridge/pci_target_unit/del_sync/N1243/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C11/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1243/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C10/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1243/FROM ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C11/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/del_sync/N1243/LOGIC_ZERO_260 (
      .O (\bridge/pci_target_unit/del_sync/N1243/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1243/YUSED (
      .I (\bridge/pci_target_unit/del_sync/N1243/XORG ),
      .O (\bridge/pci_target_unit/del_sync/N1244 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1243/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1243/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1243 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1243/COUTUSED (
      .I (\bridge/pci_target_unit/del_sync/N1243/CYMUXG ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C12/C1/O )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<2> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [2])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<3> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [3])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[3]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[3]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C14/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C13/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1245/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1245/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C14/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1245/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C13/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1245/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1245/CYMUXG )
    );
    defparam \bridge/pci_target_unit/del_sync/N1245/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1245/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_cycle_count [11]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1245/GROM )
    );
    defparam \bridge/pci_target_unit/del_sync/N1245/F .INIT = 16'hFF00;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1245/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/comp_cycle_count [10]),
      .O (\bridge/pci_target_unit/del_sync/N1245/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C13/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C12/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1245/FROM ),
      .O (\bridge/pci_target_unit/del_sync/N1245/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C13/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1245/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C12/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1245/FROM ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C13/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/del_sync/N1245/LOGIC_ZERO_261 (
      .O (\bridge/pci_target_unit/del_sync/N1245/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1245/YUSED (
      .I (\bridge/pci_target_unit/del_sync/N1245/XORG ),
      .O (\bridge/pci_target_unit/del_sync/N1246 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1245/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1245/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1245 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1245/COUTUSED (
      .I (\bridge/pci_target_unit/del_sync/N1245/CYMUXG ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C14/C1/O )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_outTransactionCount<0>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/SRNOT )
    );
    X_INV \bridge/pci_target_unit/fifos/pciw_outTransactionCount<0>/BYMUX (
      .I (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [0]),
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/BYNOT )
    );
    X_FF \bridge/pci_target_unit/fifos/pciw_outTransactionCount_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/BYNOT ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/FFY/ASYNC_FF_GSR_OR )
      ,
      .O (\bridge/pci_target_unit/fifos/pciw_outTransactionCount [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pciw_outTransactionCount<0>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pciw_outTransactionCount[0]/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C16/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C15/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1247/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1247/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C16/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1247/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C15/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1247/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1247/CYMUXG )
    );
    defparam \bridge/pci_target_unit/del_sync/N1247/G .INIT = 16'hCCCC;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1247/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/comp_cycle_count [13]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1247/GROM )
    );
    defparam \bridge/pci_target_unit/del_sync/N1247/F .INIT = 16'hFF00;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1247/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/del_sync/comp_cycle_count [12]),
      .O (\bridge/pci_target_unit/del_sync/N1247/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C15/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C14/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1247/FROM ),
      .O (\bridge/pci_target_unit/del_sync/N1247/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C15/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1247/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C14/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1247/FROM ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C15/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/del_sync/N1247/LOGIC_ZERO_262 (
      .O (\bridge/pci_target_unit/del_sync/N1247/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1247/YUSED (
      .I (\bridge/pci_target_unit/del_sync/N1247/XORG ),
      .O (\bridge/pci_target_unit/del_sync/N1248 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1247/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1247/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1247 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1247/COUTUSED (
      .I (\bridge/pci_target_unit/del_sync/N1247/CYMUXG ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C16/C1/O )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C18/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C17/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1249/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1249/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C18/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1249/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C17/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1249/GROM ),
      .O (\bridge/pci_target_unit/del_sync/N1249/CYMUXG )
    );
    defparam \bridge/pci_target_unit/del_sync/N1249/G .INIT = 16'hF0F0;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1249/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_cycle_count [15]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1249/GROM )
    );
    defparam \bridge/pci_target_unit/del_sync/N1249/F .INIT = 16'hCCCC;
    X_LUT4 \bridge/pci_target_unit/del_sync/N1249/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/del_sync/comp_cycle_count [14]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/N1249/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C17/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C16/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/N1249/FROM ),
      .O (\bridge/pci_target_unit/del_sync/N1249/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/del_sync/C1264/C17/C1 (
      .IA (\bridge/pci_target_unit/del_sync/N1249/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/del_sync/C1264/C16/C1/O ),
      .SEL (\bridge/pci_target_unit/del_sync/N1249/FROM ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C17/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/del_sync/N1249/LOGIC_ZERO_263 (
      .O (\bridge/pci_target_unit/del_sync/N1249/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1249/YUSED (
      .I (\bridge/pci_target_unit/del_sync/N1249/XORG ),
      .O (\bridge/pci_target_unit/del_sync/N1250 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1249/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1249/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1249 )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1249/COUTUSED (
      .I (\bridge/pci_target_unit/del_sync/N1249/CYMUXG ),
      .O (\bridge/pci_target_unit/del_sync/C1264/C18/C1/O )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[5]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<4> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [4])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<5> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [5]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [5])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[5]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/pci_target_unit/del_sync/comp_cycle_count<16>_rt .INIT = 16'hF0F0;
    X_LUT4 \bridge/pci_target_unit/del_sync/comp_cycle_count<16>_rt (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/del_sync/comp_cycle_count [16]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/del_sync/comp_cycle_count[16]_rt )
    );
    X_XOR2 \bridge/pci_target_unit/del_sync/C1264/C19/C0 (
      .I0 (\bridge/pci_target_unit/del_sync/C1264/C18/C1/O ),
      .I1 (\bridge/pci_target_unit/del_sync/comp_cycle_count[16]_rt ),
      .O (\bridge/pci_target_unit/del_sync/N1251/XORF )
    );
    X_BUF \bridge/pci_target_unit/del_sync/N1251/XUSED (
      .I (\bridge/pci_target_unit/del_sync/N1251/XORF ),
      .O (\bridge/pci_target_unit/del_sync/N1251 )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C4/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C3/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1717/GROM ),
      .O (\CRT/ssvga_wbm_if/N1717/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C4/C1 (
      .IA (\CRT/ssvga_wbm_if/N1717/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C3/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1717/GROM ),
      .O (\CRT/ssvga_wbm_if/N1717/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1717/G .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_wbm_if/N1717/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [3]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1717/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1717/F .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_wbm_if/N1717/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [2]),
      .O (\CRT/ssvga_wbm_if/N1717/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C3/C0 (
      .I0 (\CRT/ssvga_wbm_if/N1717/LOGIC_ONE ),
      .I1 (\CRT/ssvga_wbm_if/N1717/FROM ),
      .O (\CRT/ssvga_wbm_if/N1717/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C3/C1 (
      .IA (\CRT/ssvga_wbm_if/N1717/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/N1717/LOGIC_ONE ),
      .SEL (\CRT/ssvga_wbm_if/N1717/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C3/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1717/LOGIC_ZERO_264 (
      .O (\CRT/ssvga_wbm_if/N1717/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1717/YUSED (
      .I (\CRT/ssvga_wbm_if/N1717/XORG ),
      .O (\CRT/ssvga_wbm_if/N1718 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1717/XUSED (
      .I (\CRT/ssvga_wbm_if/N1717/XORF ),
      .O (\CRT/ssvga_wbm_if/N1717 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1717/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1717/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C4/C1/O )
    );
    X_ONE \CRT/ssvga_wbm_if/N1717/LOGIC_ONE_265 (
      .O (\CRT/ssvga_wbm_if/N1717/LOGIC_ONE )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C6/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C5/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1719/GROM ),
      .O (\CRT/ssvga_wbm_if/N1719/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C6/C1 (
      .IA (\CRT/ssvga_wbm_if/N1719/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C5/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1719/GROM ),
      .O (\CRT/ssvga_wbm_if/N1719/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1719/G .INIT = 16'hAAAA;
    X_LUT4 \CRT/ssvga_wbm_if/N1719/G (
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1719/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1719/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_wbm_if/N1719/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [4]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1719/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C5/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C4/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1719/FROM ),
      .O (\CRT/ssvga_wbm_if/N1719/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C5/C1 (
      .IA (\CRT/ssvga_wbm_if/N1719/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C4/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1719/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C5/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1719/LOGIC_ZERO_266 (
      .O (\CRT/ssvga_wbm_if/N1719/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1719/YUSED (
      .I (\CRT/ssvga_wbm_if/N1719/XORG ),
      .O (\CRT/ssvga_wbm_if/N1720 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1719/XUSED (
      .I (\CRT/ssvga_wbm_if/N1719/XORF ),
      .O (\CRT/ssvga_wbm_if/N1719 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1719/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1719/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C6/C1/O )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[7]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<6> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [6])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<7> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [7]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [7])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[7]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[7]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C8/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C7/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1721/GROM ),
      .O (\CRT/ssvga_wbm_if/N1721/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C8/C1 (
      .IA (\CRT/ssvga_wbm_if/N1721/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C7/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1721/GROM ),
      .O (\CRT/ssvga_wbm_if/N1721/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1721/G .INIT = 16'hAAAA;
    X_LUT4 \CRT/ssvga_wbm_if/N1721/G (
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1721/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1721/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1721/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [6]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1721/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C7/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C6/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1721/FROM ),
      .O (\CRT/ssvga_wbm_if/N1721/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C7/C1 (
      .IA (\CRT/ssvga_wbm_if/N1721/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C6/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1721/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C7/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1721/LOGIC_ZERO_267 (
      .O (\CRT/ssvga_wbm_if/N1721/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1721/YUSED (
      .I (\CRT/ssvga_wbm_if/N1721/XORG ),
      .O (\CRT/ssvga_wbm_if/N1722 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1721/XUSED (
      .I (\CRT/ssvga_wbm_if/N1721/XORF ),
      .O (\CRT/ssvga_wbm_if/N1721 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1721/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1721/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C8/C1/O )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C10/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C9/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1723/GROM ),
      .O (\CRT/ssvga_wbm_if/N1723/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C10/C1 (
      .IA (\CRT/ssvga_wbm_if/N1723/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C9/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1723/GROM ),
      .O (\CRT/ssvga_wbm_if/N1723/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1723/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1723/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [9]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1723/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1723/F .INIT = 16'hAAAA;
    X_LUT4 \CRT/ssvga_wbm_if/N1723/F (
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [8]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1723/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C9/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C8/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1723/FROM ),
      .O (\CRT/ssvga_wbm_if/N1723/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C9/C1 (
      .IA (\CRT/ssvga_wbm_if/N1723/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C8/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1723/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C9/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1723/LOGIC_ZERO_268 (
      .O (\CRT/ssvga_wbm_if/N1723/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1723/YUSED (
      .I (\CRT/ssvga_wbm_if/N1723/XORG ),
      .O (\CRT/ssvga_wbm_if/N1724 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1723/XUSED (
      .I (\CRT/ssvga_wbm_if/N1723/XORF ),
      .O (\CRT/ssvga_wbm_if/N1723 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1723/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1723/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C10/C1/O )
    );
    X_INV \bridge/pci_target_unit/pcit_if_addr_out<9>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[9]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<8> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[9]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [8])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<9>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[9]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/pci_target_if/norm_address_reg<9> (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [9]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/pcit_sm_addr_phase_out ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/pcit_if_addr_out[9]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/pcit_if_addr_out [9])
    );
    X_OR2 \bridge/pci_target_unit/pcit_if_addr_out<9>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/pcit_if_addr_out[9]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/pcit_if_addr_out[9]/FFX/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C12/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C11/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1725/GROM ),
      .O (\CRT/ssvga_wbm_if/N1725/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C12/C1 (
      .IA (\CRT/ssvga_wbm_if/N1725/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C11/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1725/GROM ),
      .O (\CRT/ssvga_wbm_if/N1725/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1725/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_wbm_if/N1725/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [11]),
      .O (\CRT/ssvga_wbm_if/N1725/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1725/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1725/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [10]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1725/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C11/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C10/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1725/FROM ),
      .O (\CRT/ssvga_wbm_if/N1725/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C11/C1 (
      .IA (\CRT/ssvga_wbm_if/N1725/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C10/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1725/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C11/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1725/LOGIC_ZERO_269 (
      .O (\CRT/ssvga_wbm_if/N1725/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1725/YUSED (
      .I (\CRT/ssvga_wbm_if/N1725/XORG ),
      .O (\CRT/ssvga_wbm_if/N1726 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1725/XUSED (
      .I (\CRT/ssvga_wbm_if/N1725/XORF ),
      .O (\CRT/ssvga_wbm_if/N1725 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1725/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1725/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C12/C1/O )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C14/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C13/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1727/GROM ),
      .O (\CRT/ssvga_wbm_if/N1727/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C14/C1 (
      .IA (\CRT/ssvga_wbm_if/N1727/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C13/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1727/GROM ),
      .O (\CRT/ssvga_wbm_if/N1727/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1727/G .INIT = 16'hAAAA;
    X_LUT4 \CRT/ssvga_wbm_if/N1727/G (
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [13]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1727/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1727/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_wbm_if/N1727/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [12]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1727/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C13/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C12/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1727/FROM ),
      .O (\CRT/ssvga_wbm_if/N1727/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C13/C1 (
      .IA (\CRT/ssvga_wbm_if/N1727/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C12/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1727/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C13/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1727/LOGIC_ZERO_270 (
      .O (\CRT/ssvga_wbm_if/N1727/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1727/YUSED (
      .I (\CRT/ssvga_wbm_if/N1727/XORG ),
      .O (\CRT/ssvga_wbm_if/N1728 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1727/XUSED (
      .I (\CRT/ssvga_wbm_if/N1727/XORF ),
      .O (\CRT/ssvga_wbm_if/N1727 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1727/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1727/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C14/C1/O )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<4>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[4]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next_reg<4> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_waddr [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wallow ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next [4])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[4]/SRNOT )
      ,
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wgrey_next[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C16/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C15/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1729/GROM ),
      .O (\CRT/ssvga_wbm_if/N1729/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C16/C1 (
      .IA (\CRT/ssvga_wbm_if/N1729/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C15/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1729/GROM ),
      .O (\CRT/ssvga_wbm_if/N1729/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1729/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1729/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [15]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1729/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1729/F .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_wbm_if/N1729/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [14]),
      .O (\CRT/ssvga_wbm_if/N1729/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C15/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C14/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1729/FROM ),
      .O (\CRT/ssvga_wbm_if/N1729/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C15/C1 (
      .IA (\CRT/ssvga_wbm_if/N1729/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C14/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1729/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C15/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1729/LOGIC_ZERO_271 (
      .O (\CRT/ssvga_wbm_if/N1729/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1729/YUSED (
      .I (\CRT/ssvga_wbm_if/N1729/XORG ),
      .O (\CRT/ssvga_wbm_if/N1730 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1729/XUSED (
      .I (\CRT/ssvga_wbm_if/N1729/XORF ),
      .O (\CRT/ssvga_wbm_if/N1729 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1729/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1729/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C16/C1/O )
    );
    X_INV \bridge/out_bckp_irdy_en_out/SRMUX (
      .I (N_RST),
      .O (\bridge/out_bckp_irdy_en_out/SRNOT )
    );
    X_FF \bridge/output_backup/irdy_en_out_reg (
      .I (\bridge/out_bckp_frame_en_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/out_bckp_irdy_en_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/out_bckp_irdy_en_out )
    );
    X_OR2 \bridge/out_bckp_irdy_en_out/FFY/ASYNC_FF_GSR_OR_272 (
      .I0 (\bridge/out_bckp_irdy_en_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/out_bckp_irdy_en_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C18/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C17/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1731/GROM ),
      .O (\CRT/ssvga_wbm_if/N1731/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C18/C1 (
      .IA (\CRT/ssvga_wbm_if/N1731/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C17/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1731/GROM ),
      .O (\CRT/ssvga_wbm_if/N1731/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1731/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1731/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [17]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1731/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1731/F .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_wbm_if/N1731/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [16]),
      .O (\CRT/ssvga_wbm_if/N1731/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C17/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C16/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1731/FROM ),
      .O (\CRT/ssvga_wbm_if/N1731/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C17/C1 (
      .IA (\CRT/ssvga_wbm_if/N1731/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C16/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1731/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C17/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1731/LOGIC_ZERO_273 (
      .O (\CRT/ssvga_wbm_if/N1731/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1731/YUSED (
      .I (\CRT/ssvga_wbm_if/N1731/XORG ),
      .O (\CRT/ssvga_wbm_if/N1732 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1731/XUSED (
      .I (\CRT/ssvga_wbm_if/N1731/XORF ),
      .O (\CRT/ssvga_wbm_if/N1731 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1731/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1731/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C18/C1/O )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C20/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C19/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1733/GROM ),
      .O (\CRT/ssvga_wbm_if/N1733/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C20/C1 (
      .IA (\CRT/ssvga_wbm_if/N1733/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C19/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1733/GROM ),
      .O (\CRT/ssvga_wbm_if/N1733/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1733/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1733/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [19]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1733/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1733/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1733/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [18]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1733/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C19/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C18/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1733/FROM ),
      .O (\CRT/ssvga_wbm_if/N1733/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C19/C1 (
      .IA (\CRT/ssvga_wbm_if/N1733/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C18/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1733/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C19/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1733/LOGIC_ZERO_274 (
      .O (\CRT/ssvga_wbm_if/N1733/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1733/YUSED (
      .I (\CRT/ssvga_wbm_if/N1733/XORG ),
      .O (\CRT/ssvga_wbm_if/N1734 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1733/XUSED (
      .I (\CRT/ssvga_wbm_if/N1733/XORF ),
      .O (\CRT/ssvga_wbm_if/N1733 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1733/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1733/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C20/C1/O )
    );
    X_INV \bridge/parity_checker/check_perr/SRMUX (
      .I (N_RST),
      .O (\bridge/parity_checker/check_perr/SRNOT )
    );
    X_FF \bridge/parity_checker/check_perr_reg (
      .I (\bridge/out_bckp_par_en_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST (\bridge/parity_checker/check_perr/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/parity_checker/check_perr )
    );
    X_OR2 \bridge/parity_checker/check_perr/FFY/ASYNC_FF_GSR_OR_275 (
      .I0 (\bridge/parity_checker/check_perr/SRNOT ),
      .I1 (GSR),
      .O (\bridge/parity_checker/check_perr/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C22/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C21/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1735/GROM ),
      .O (\CRT/ssvga_wbm_if/N1735/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C22/C1 (
      .IA (\CRT/ssvga_wbm_if/N1735/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C21/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1735/GROM ),
      .O (\CRT/ssvga_wbm_if/N1735/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1735/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1735/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [21]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1735/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1735/F .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_wbm_if/N1735/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [20]),
      .O (\CRT/ssvga_wbm_if/N1735/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C21/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C20/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1735/FROM ),
      .O (\CRT/ssvga_wbm_if/N1735/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C21/C1 (
      .IA (\CRT/ssvga_wbm_if/N1735/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C20/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1735/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C21/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1735/LOGIC_ZERO_276 (
      .O (\CRT/ssvga_wbm_if/N1735/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1735/YUSED (
      .I (\CRT/ssvga_wbm_if/N1735/XORG ),
      .O (\CRT/ssvga_wbm_if/N1736 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1735/XUSED (
      .I (\CRT/ssvga_wbm_if/N1735/XORF ),
      .O (\CRT/ssvga_wbm_if/N1735 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1735/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1735/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C22/C1/O )
    );
    X_INV \bridge/pci_target_unit/del_sync/sync_comp_req_pending/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/sync_comp_req_pending/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/req_sync/sync_data_out_reg<0> (
      .I (\bridge/pci_target_unit/pcit_if_read_processing_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/sync_comp_req_pending/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/sync_comp_req_pending )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/sync_comp_req_pending/FFY/ASYNC_FF_GSR_OR_277 (
      .I0 (\bridge/pci_target_unit/del_sync/sync_comp_req_pending/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/sync_comp_req_pending/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C24/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C23/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1737/GROM ),
      .O (\CRT/ssvga_wbm_if/N1737/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C24/C1 (
      .IA (\CRT/ssvga_wbm_if/N1737/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C23/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1737/GROM ),
      .O (\CRT/ssvga_wbm_if/N1737/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1737/G .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_wbm_if/N1737/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [23]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1737/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1737/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1737/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [22]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1737/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C23/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C22/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1737/FROM ),
      .O (\CRT/ssvga_wbm_if/N1737/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C23/C1 (
      .IA (\CRT/ssvga_wbm_if/N1737/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C22/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1737/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C23/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1737/LOGIC_ZERO_278 (
      .O (\CRT/ssvga_wbm_if/N1737/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1737/YUSED (
      .I (\CRT/ssvga_wbm_if/N1737/XORG ),
      .O (\CRT/ssvga_wbm_if/N1738 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1737/XUSED (
      .I (\CRT/ssvga_wbm_if/N1737/XORF ),
      .O (\CRT/ssvga_wbm_if/N1737 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1737/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1737/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C24/C1/O )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/req_sync/sync_data_out_reg<0> (
      .I (\bridge/wishbone_slave_unit/del_sync_req_req_pending_out ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending/FFY/ASYNC_FF_GSR_OR_279 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync/sync_comp_req_pending/FFY/ASYNC_FF_GSR_OR )

    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C26/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C25/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1739/GROM ),
      .O (\CRT/ssvga_wbm_if/N1739/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C26/C1 (
      .IA (\CRT/ssvga_wbm_if/N1739/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C25/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1739/GROM ),
      .O (\CRT/ssvga_wbm_if/N1739/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1739/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_wbm_if/N1739/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [25]),
      .O (\CRT/ssvga_wbm_if/N1739/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1739/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1739/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [24]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1739/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C25/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C24/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1739/FROM ),
      .O (\CRT/ssvga_wbm_if/N1739/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C25/C1 (
      .IA (\CRT/ssvga_wbm_if/N1739/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C24/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1739/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C25/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1739/LOGIC_ZERO_280 (
      .O (\CRT/ssvga_wbm_if/N1739/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1739/YUSED (
      .I (\CRT/ssvga_wbm_if/N1739/XORG ),
      .O (\CRT/ssvga_wbm_if/N1740 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1739/XUSED (
      .I (\CRT/ssvga_wbm_if/N1739/XORF ),
      .O (\CRT/ssvga_wbm_if/N1739 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1739/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1739/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C26/C1/O )
    );
    X_INV \crt_vsync/SRMUX (
      .I (N_RST),
      .O (\crt_vsync/SRNOT )
    );
    X_INV \crt_vsync/BYMUX (
      .I (\CRT/ssvga_crtc/vcntr [2]),
      .O (\crt_vsync/BYNOT )
    );
    X_FF \CRT/ssvga_crtc/vsync_reg (
      .I (\crt_vsync/BYNOT ),
      .CLK (CRT_CLK_BUFGPed),
      .CE (N12163),
      .SET (GND),
      .RST (\crt_vsync/FFY/ASYNC_FF_GSR_OR ),
      .O (crt_vsync)
    );
    X_OR2 \crt_vsync/FFY/ASYNC_FF_GSR_OR_281 (
      .I0 (\crt_vsync/SRNOT ),
      .I1 (GSR),
      .O (\crt_vsync/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C28/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C27/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1741/GROM ),
      .O (\CRT/ssvga_wbm_if/N1741/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C28/C1 (
      .IA (\CRT/ssvga_wbm_if/N1741/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C27/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1741/GROM ),
      .O (\CRT/ssvga_wbm_if/N1741/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1741/G .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_wbm_if/N1741/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [27]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1741/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1741/F .INIT = 16'hAAAA;
    X_LUT4 \CRT/ssvga_wbm_if/N1741/F (
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [26]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1741/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C27/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C26/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1741/FROM ),
      .O (\CRT/ssvga_wbm_if/N1741/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C27/C1 (
      .IA (\CRT/ssvga_wbm_if/N1741/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C26/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1741/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C27/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1741/LOGIC_ZERO_282 (
      .O (\CRT/ssvga_wbm_if/N1741/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1741/YUSED (
      .I (\CRT/ssvga_wbm_if/N1741/XORG ),
      .O (\CRT/ssvga_wbm_if/N1742 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1741/XUSED (
      .I (\CRT/ssvga_wbm_if/N1741/XORF ),
      .O (\CRT/ssvga_wbm_if/N1741 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1741/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1741/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C28/C1/O )
    );
    X_INV \bridge/conf_perr_response_out/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_perr_response_out/SRNOT )
    );
    X_FF \bridge/configuration/command_bit6_reg (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [6]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C281/N3 ),
      .SET (GND),
      .RST (\bridge/conf_perr_response_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_perr_response_out )
    );
    X_OR2 \bridge/conf_perr_response_out/FFY/ASYNC_FF_GSR_OR_283 (
      .I0 (\bridge/conf_perr_response_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_perr_response_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C30/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C29/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1743/GROM ),
      .O (\CRT/ssvga_wbm_if/N1743/XORG )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C30/C1 (
      .IA (\CRT/ssvga_wbm_if/N1743/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C29/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1743/GROM ),
      .O (\CRT/ssvga_wbm_if/N1743/CYMUXG )
    );
    defparam \CRT/ssvga_wbm_if/N1743/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_wbm_if/N1743/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [29]),
      .O (\CRT/ssvga_wbm_if/N1743/GROM )
    );
    defparam \CRT/ssvga_wbm_if/N1743/F .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_wbm_if/N1743/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [28]),
      .O (\CRT/ssvga_wbm_if/N1743/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C29/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C28/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1743/FROM ),
      .O (\CRT/ssvga_wbm_if/N1743/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C29/C1 (
      .IA (\CRT/ssvga_wbm_if/N1743/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C28/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1743/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C29/C1/O )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1743/LOGIC_ZERO_284 (
      .O (\CRT/ssvga_wbm_if/N1743/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_wbm_if/N1743/YUSED (
      .I (\CRT/ssvga_wbm_if/N1743/XORG ),
      .O (\CRT/ssvga_wbm_if/N1744 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1743/XUSED (
      .I (\CRT/ssvga_wbm_if/N1743/XORF ),
      .O (\CRT/ssvga_wbm_if/N1743 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1743/COUTUSED (
      .I (\CRT/ssvga_wbm_if/N1743/CYMUXG ),
      .O (\CRT/ssvga_wbm_if/C1473/C30/C1/O )
    );
    X_INV \bridge/pci_target_unit/del_sync/comp_done_reg_main/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/del_sync/comp_done_reg_main/SRNOT )
    );
    X_FF \bridge/pci_target_unit/del_sync/comp_done_reg_main_reg (
      .I (\bridge/pci_target_unit/del_sync/sync_comp_done ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/del_sync/comp_done_reg_main/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/del_sync/comp_done_reg_main )
    );
    X_OR2
     \bridge/pci_target_unit/del_sync/comp_done_reg_main/FFY/ASYNC_FF_GSR_OR_285 (
      .I0 (\bridge/pci_target_unit/del_sync/comp_done_reg_main/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/del_sync/comp_done_reg_main/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C32/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C31/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]_rt ),
      .O (\CRT/ssvga_wbm_if/N1745/XORG )
    );
    defparam \bridge/wishbone_slave_unit/wb_addr_dec/addr1<31>_rt .INIT = 16'hAAAA;
    X_LUT4 \bridge/wishbone_slave_unit/wb_addr_dec/addr1<31>_rt (
      .ADR0 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [31]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/wb_addr_dec/addr1[31]_rt )
    );
    defparam \CRT/ssvga_wbm_if/N1745/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_wbm_if/N1745/F (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/wb_addr_dec/addr1 [30]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_wbm_if/N1745/FROM )
    );
    X_XOR2 \CRT/ssvga_wbm_if/C1473/C31/C0 (
      .I0 (\CRT/ssvga_wbm_if/C1473/C30/C1/O ),
      .I1 (\CRT/ssvga_wbm_if/N1745/FROM ),
      .O (\CRT/ssvga_wbm_if/N1745/XORF )
    );
    X_MUX2 \CRT/ssvga_wbm_if/C1473/C31/C1 (
      .IA (\CRT/ssvga_wbm_if/N1745/LOGIC_ZERO ),
      .IB (\CRT/ssvga_wbm_if/C1473/C30/C1/O ),
      .SEL (\CRT/ssvga_wbm_if/N1745/FROM ),
      .O (\CRT/ssvga_wbm_if/C1473/C31/C1/O )
    );
    X_BUF \CRT/ssvga_wbm_if/N1745/YUSED (
      .I (\CRT/ssvga_wbm_if/N1745/XORG ),
      .O (\CRT/ssvga_wbm_if/N1746 )
    );
    X_BUF \CRT/ssvga_wbm_if/N1745/XUSED (
      .I (\CRT/ssvga_wbm_if/N1745/XORF ),
      .O (\CRT/ssvga_wbm_if/N1745 )
    );
    X_ZERO \CRT/ssvga_wbm_if/N1745/LOGIC_ZERO_286 (
      .O (\CRT/ssvga_wbm_if/N1745/LOGIC_ZERO )
    );
    X_XOR2 \CRT/ssvga_crtc/C529/C4/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C3/C1/O ),
      .I1 (\CRT/ssvga_crtc/N326/GROM ),
      .O (\CRT/ssvga_crtc/N326/XORG )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C4/C1 (
      .IA (\CRT/ssvga_crtc/N326/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C529/C3/C1/O ),
      .SEL (\CRT/ssvga_crtc/N326/GROM ),
      .O (\CRT/ssvga_crtc/N326/CYMUXG )
    );
    defparam \CRT/ssvga_crtc/N326/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_crtc/N326/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/vcntr [1]),
      .O (\CRT/ssvga_crtc/N326/GROM )
    );
    defparam \CRT/ssvga_crtc/N326/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_crtc/N326/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/vcntr [0]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N326/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C529/C3/C0 (
      .I0 (\CRT/ssvga_crtc/N326/LOGIC_ONE ),
      .I1 (\CRT/ssvga_crtc/N326/FROM ),
      .O (\CRT/ssvga_crtc/N326/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C3/C1 (
      .IA (\CRT/ssvga_crtc/N326/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/N326/LOGIC_ONE ),
      .SEL (\CRT/ssvga_crtc/N326/FROM ),
      .O (\CRT/ssvga_crtc/C529/C3/C1/O )
    );
    X_ZERO \CRT/ssvga_crtc/N326/LOGIC_ZERO_287 (
      .O (\CRT/ssvga_crtc/N326/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_crtc/N326/YUSED (
      .I (\CRT/ssvga_crtc/N326/XORG ),
      .O (\CRT/ssvga_crtc/N327 )
    );
    X_BUF \CRT/ssvga_crtc/N326/XUSED (
      .I (\CRT/ssvga_crtc/N326/XORF ),
      .O (\CRT/ssvga_crtc/N326 )
    );
    X_BUF \CRT/ssvga_crtc/N326/COUTUSED (
      .I (\CRT/ssvga_crtc/N326/CYMUXG ),
      .O (\CRT/ssvga_crtc/C529/C4/C1/O )
    );
    X_ONE \CRT/ssvga_crtc/N326/LOGIC_ONE_288 (
      .O (\CRT/ssvga_crtc/N326/LOGIC_ONE )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [0])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[1]/FFX/ASYNC_FF_GSR_OR )

    );
    X_XOR2 \CRT/ssvga_crtc/C529/C6/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C5/C1/O ),
      .I1 (\CRT/ssvga_crtc/N328/GROM ),
      .O (\CRT/ssvga_crtc/N328/XORG )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C6/C1 (
      .IA (\CRT/ssvga_crtc/N328/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C529/C5/C1/O ),
      .SEL (\CRT/ssvga_crtc/N328/GROM ),
      .O (\CRT/ssvga_crtc/N328/CYMUXG )
    );
    defparam \CRT/ssvga_crtc/N328/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_crtc/N328/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/vcntr [3]),
      .O (\CRT/ssvga_crtc/N328/GROM )
    );
    defparam \CRT/ssvga_crtc/N328/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_crtc/N328/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/vcntr [2]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N328/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C529/C5/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C4/C1/O ),
      .I1 (\CRT/ssvga_crtc/N328/FROM ),
      .O (\CRT/ssvga_crtc/N328/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C5/C1 (
      .IA (\CRT/ssvga_crtc/N328/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C529/C4/C1/O ),
      .SEL (\CRT/ssvga_crtc/N328/FROM ),
      .O (\CRT/ssvga_crtc/C529/C5/C1/O )
    );
    X_ZERO \CRT/ssvga_crtc/N328/LOGIC_ZERO_289 (
      .O (\CRT/ssvga_crtc/N328/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_crtc/N328/YUSED (
      .I (\CRT/ssvga_crtc/N328/XORG ),
      .O (\CRT/ssvga_crtc/N329 )
    );
    X_BUF \CRT/ssvga_crtc/N328/XUSED (
      .I (\CRT/ssvga_crtc/N328/XORF ),
      .O (\CRT/ssvga_crtc/N328 )
    );
    X_BUF \CRT/ssvga_crtc/N328/COUTUSED (
      .I (\CRT/ssvga_crtc/N328/CYMUXG ),
      .O (\CRT/ssvga_crtc/C529/C6/C1/O )
    );
    X_XOR2 \CRT/ssvga_crtc/C529/C8/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C7/C1/O ),
      .I1 (\CRT/ssvga_crtc/N330/GROM ),
      .O (\CRT/ssvga_crtc/N330/XORG )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C8/C1 (
      .IA (\CRT/ssvga_crtc/N330/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C529/C7/C1/O ),
      .SEL (\CRT/ssvga_crtc/N330/GROM ),
      .O (\CRT/ssvga_crtc/N330/CYMUXG )
    );
    defparam \CRT/ssvga_crtc/N330/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_crtc/N330/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/vcntr [5]),
      .O (\CRT/ssvga_crtc/N330/GROM )
    );
    defparam \CRT/ssvga_crtc/N330/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_crtc/N330/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/vcntr [4]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N330/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C529/C7/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C6/C1/O ),
      .I1 (\CRT/ssvga_crtc/N330/FROM ),
      .O (\CRT/ssvga_crtc/N330/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C7/C1 (
      .IA (\CRT/ssvga_crtc/N330/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C529/C6/C1/O ),
      .SEL (\CRT/ssvga_crtc/N330/FROM ),
      .O (\CRT/ssvga_crtc/C529/C7/C1/O )
    );
    X_ZERO \CRT/ssvga_crtc/N330/LOGIC_ZERO_290 (
      .O (\CRT/ssvga_crtc/N330/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_crtc/N330/YUSED (
      .I (\CRT/ssvga_crtc/N330/XORG ),
      .O (\CRT/ssvga_crtc/N331 )
    );
    X_BUF \CRT/ssvga_crtc/N330/XUSED (
      .I (\CRT/ssvga_crtc/N330/XORF ),
      .O (\CRT/ssvga_crtc/N330 )
    );
    X_BUF \CRT/ssvga_crtc/N330/COUTUSED (
      .I (\CRT/ssvga_crtc/N330/CYMUXG ),
      .O (\CRT/ssvga_crtc/C529/C8/C1/O )
    );
    defparam \bridge/pci_io_mux/ad_en_low_gen/C0 .INIT = 16'h0505;
    X_LUT4 \bridge/pci_io_mux/ad_en_low_gen/C0 (
      .ADR0 (\bridge/pci_mux_tar_ad_en_in ),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_mux_mas_ad_en_in ),
      .ADR3 (VCC),
      .O (\N12322/GROM )
    );
    defparam \bridge/pci_io_mux/ad_en_mlow_gen/C0 .INIT = 16'h0055;
    X_LUT4 \bridge/pci_io_mux/ad_en_mlow_gen/C0 (
      .ADR0 (\bridge/pci_mux_tar_ad_en_in ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_mux_mas_ad_en_in ),
      .O (\N12322/FROM )
    );
    X_BUF \N12322/YUSED (
      .I (\N12322/GROM ),
      .O (N12314)
    );
    X_BUF \N12322/XUSED (
      .I (\N12322/FROM ),
      .O (N12322)
    );
    X_XOR2 \CRT/ssvga_crtc/C529/C10/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C9/C1/O ),
      .I1 (\CRT/ssvga_crtc/N332/GROM ),
      .O (\CRT/ssvga_crtc/N332/XORG )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C10/C1 (
      .IA (\CRT/ssvga_crtc/N332/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C529/C9/C1/O ),
      .SEL (\CRT/ssvga_crtc/N332/GROM ),
      .O (\CRT/ssvga_crtc/N332/CYMUXG )
    );
    defparam \CRT/ssvga_crtc/N332/G .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_crtc/N332/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/vcntr [7]),
      .O (\CRT/ssvga_crtc/N332/GROM )
    );
    defparam \CRT/ssvga_crtc/N332/F .INIT = 16'hAAAA;
    X_LUT4 \CRT/ssvga_crtc/N332/F (
      .ADR0 (\CRT/ssvga_crtc/vcntr [6]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N332/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C529/C9/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C8/C1/O ),
      .I1 (\CRT/ssvga_crtc/N332/FROM ),
      .O (\CRT/ssvga_crtc/N332/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C9/C1 (
      .IA (\CRT/ssvga_crtc/N332/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C529/C8/C1/O ),
      .SEL (\CRT/ssvga_crtc/N332/FROM ),
      .O (\CRT/ssvga_crtc/C529/C9/C1/O )
    );
    X_ZERO \CRT/ssvga_crtc/N332/LOGIC_ZERO_291 (
      .O (\CRT/ssvga_crtc/N332/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_crtc/N332/YUSED (
      .I (\CRT/ssvga_crtc/N332/XORG ),
      .O (\CRT/ssvga_crtc/N333 )
    );
    X_BUF \CRT/ssvga_crtc/N332/XUSED (
      .I (\CRT/ssvga_crtc/N332/XORF ),
      .O (\CRT/ssvga_crtc/N332 )
    );
    X_BUF \CRT/ssvga_crtc/N332/COUTUSED (
      .I (\CRT/ssvga_crtc/N332/CYMUXG ),
      .O (\CRT/ssvga_crtc/C529/C10/C1/O )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [2])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr<3>/FFY/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFY/RST )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [3])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr<3>/FFX/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFX/RST )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[3]/FFX/ASYNC_FF_GSR_OR )

    );
    X_XOR2 \CRT/ssvga_crtc/C529/C12/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C11/C1/O ),
      .I1 (\CRT/ssvga_crtc/vcntr[9]_rt ),
      .O (\CRT/ssvga_crtc/N334/XORG )
    );
    defparam \CRT/ssvga_crtc/vcntr<9>_rt .INIT = 16'hFF00;
    X_LUT4 \CRT/ssvga_crtc/vcntr<9>_rt (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\CRT/ssvga_crtc/vcntr [9]),
      .O (\CRT/ssvga_crtc/vcntr[9]_rt )
    );
    defparam \CRT/ssvga_crtc/N334/F .INIT = 16'hAAAA;
    X_LUT4 \CRT/ssvga_crtc/N334/F (
      .ADR0 (\CRT/ssvga_crtc/vcntr [8]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N334/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C529/C11/C0 (
      .I0 (\CRT/ssvga_crtc/C529/C10/C1/O ),
      .I1 (\CRT/ssvga_crtc/N334/FROM ),
      .O (\CRT/ssvga_crtc/N334/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C529/C11/C1 (
      .IA (\CRT/ssvga_crtc/N334/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C529/C10/C1/O ),
      .SEL (\CRT/ssvga_crtc/N334/FROM ),
      .O (\CRT/ssvga_crtc/C529/C11/C1/O )
    );
    X_BUF \CRT/ssvga_crtc/N334/YUSED (
      .I (\CRT/ssvga_crtc/N334/XORG ),
      .O (\CRT/ssvga_crtc/N335 )
    );
    X_BUF \CRT/ssvga_crtc/N334/XUSED (
      .I (\CRT/ssvga_crtc/N334/XORF ),
      .O (\CRT/ssvga_crtc/N334 )
    );
    X_ZERO \CRT/ssvga_crtc/N334/LOGIC_ZERO_292 (
      .O (\CRT/ssvga_crtc/N334/LOGIC_ZERO )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3410/C4/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3410/C3/C1/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/C3413/N12 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3068/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3410/C4/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3410/C3/C1/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/C3413/N12 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3068/CYMUXG )
    );
    defparam C19090.INIT = 16'hFFF0;
    X_LUT4 C19090(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn19555),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3069 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3413/N12 )
    );
    defparam C19091.INIT = 16'hFFAA;
    X_LUT4 C19091(
      .ADR0 (syn19555),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3068 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3413/N6 )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3410/C3/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ONE ),
      .I1 (\bridge/pci_target_unit/wishbone_master/C3413/N6 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3068/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3410/C3/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ONE ),
      .SEL (\bridge/pci_target_unit/wishbone_master/C3413/N6 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3410/C3/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ZERO_293 (
      .O (\bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3068/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3068/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3069 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3068/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3068/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3068 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3068/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3068/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3410/C4/C1/O )
    );
    X_ONE \bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ONE_294 (
      .O (\bridge/pci_target_unit/wishbone_master/N3068/LOGIC_ONE )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3410/C6/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3410/C5/C1/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/C3413/N24 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3070/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3410/C6/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/N3070/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3410/C5/C1/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/C3413/N24 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3070/CYMUXG )
    );
    defparam C19088.INIT = 16'hFFCC;
    X_LUT4 C19088(
      .ADR0 (VCC),
      .ADR1 (syn19555),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3071 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3413/N24 )
    );
    defparam C19089.INIT = 16'hFFF0;
    X_LUT4 C19089(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (syn19555),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3070 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3413/N18 )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3410/C5/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3410/C4/C1/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/C3413/N18 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3070/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3410/C5/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/N3070/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3410/C4/C1/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/C3413/N18 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3410/C5/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/wishbone_master/N3070/LOGIC_ZERO_295 (
      .O (\bridge/pci_target_unit/wishbone_master/N3070/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3070/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3070/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3071 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3070/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3070/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3070 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3070/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3070/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3410/C6/C1/O )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr_reg<4> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [4]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr [4])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr<4>/FFY/SETOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[4]/FFY/SET )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr<4>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[4]/FFY/SET ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_addr[4]/FFY/ASYNC_FF_GSR_OR )

    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3410/C8/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3410/C7/C1/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/C3413/N36 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3072/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3410/C8/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/N3072/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3410/C7/C1/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/C3413/N36 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3072/CYMUXG )
    );
    defparam C19086.INIT = 16'hFFCC;
    X_LUT4 C19086(
      .ADR0 (VCC),
      .ADR1 (syn19555),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3073 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3413/N36 )
    );
    defparam C19087.INIT = 16'hFFCC;
    X_LUT4 C19087(
      .ADR0 (VCC),
      .ADR1 (syn19555),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3072 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3413/N30 )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3410/C7/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3410/C6/C1/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/C3413/N30 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3072/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3410/C7/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/N3072/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3410/C6/C1/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/C3413/N30 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3410/C7/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/wishbone_master/N3072/LOGIC_ZERO_296 (
      .O (\bridge/pci_target_unit/wishbone_master/N3072/LOGIC_ZERO )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3072/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3072/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3073 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3072/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3072/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3072 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3072/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3072/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3410/C8/C1/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3410/C10/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3410/C9/C1/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/C3413/N48 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3074/XORG )
    );
    defparam C19084.INIT = 16'hFFF0;
    X_LUT4 C19084(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/N3075 ),
      .ADR3 (syn19555),
      .O (\bridge/pci_target_unit/wishbone_master/C3413/N48 )
    );
    defparam C19085.INIT = 16'hFFCC;
    X_LUT4 C19085(
      .ADR0 (VCC),
      .ADR1 (syn19555),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3074 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3413/N42 )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3410/C9/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3410/C8/C1/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/C3413/N42 ),
      .O (\bridge/pci_target_unit/wishbone_master/N3074/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3410/C9/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/N3074/LOGIC_ZERO ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3410/C8/C1/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/C3413/N42 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3410/C9/C1/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3074/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3074/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3075 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3074/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3074/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3074 )
    );
    X_ZERO \bridge/pci_target_unit/wishbone_master/N3074/LOGIC_ZERO_297 (
      .O (\bridge/pci_target_unit/wishbone_master/N3074/LOGIC_ZERO )
    );
    X_INV \bridge/wishbone_slave_unit/del_sync_comp_flush_out/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/del_sync_comp_flush_out/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/del_sync/comp_flush_out_reg (
      .I (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [16]),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/del_sync_comp_flush_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/del_sync_comp_flush_out )
    );
    X_OR2
     \bridge/wishbone_slave_unit/del_sync_comp_flush_out/FFY/ASYNC_FF_GSR_OR_298 (
      .I0 (\bridge/wishbone_slave_unit/del_sync_comp_flush_out/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/del_sync_comp_flush_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C3/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C2/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2983/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2983/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C3/C2 (
      .IA (\bridge/pciu_err_addr_out[1] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C2/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2983/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2983/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2983/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2983/G (
      .ADR0 (\bridge/pciu_err_addr_out[1] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2983/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2983/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2983/F (
      .ADR0 (\bridge/pciu_err_addr_out[0] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2983/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C2/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/N2983/LOGIC_ZERO ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2983/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2983/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C2/C2 (
      .IA (\bridge/pciu_err_addr_out[0] ),
      .IB (\bridge/pci_target_unit/wishbone_master/N2983/LOGIC_ZERO ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2983/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C2/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2983/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2983/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N2984 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2983/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2983/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2983 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2983/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2983/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C3/C2/O )
    );
    X_ZERO \bridge/pci_target_unit/wishbone_master/N2983/LOGIC_ZERO_299 (
      .O (\bridge/pci_target_unit/wishbone_master/N2983/LOGIC_ZERO )
    );
    X_INV \bridge/conf_serr_enable_out/SRMUX (
      .I (N_RST),
      .O (\bridge/conf_serr_enable_out/SRNOT )
    );
    X_FF \bridge/configuration/command_bit8_reg (
      .I (\bridge/pci_target_unit/pci_target_if/address1_in [8]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/configuration/C280/N3 ),
      .SET (GND),
      .RST (\bridge/conf_serr_enable_out/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/conf_serr_enable_out )
    );
    X_OR2 \bridge/conf_serr_enable_out/FFY/ASYNC_FF_GSR_OR_300 (
      .I0 (\bridge/conf_serr_enable_out/SRNOT ),
      .I1 (GSR),
      .O (\bridge/conf_serr_enable_out/FFY/ASYNC_FF_GSR_OR )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C5/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C4/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2985/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2985/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C5/C2 (
      .IA (ADR_O[3]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C4/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2985/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2985/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2985/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2985/G (
      .ADR0 (ADR_O[3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2985/GROM )
    );
    defparam C19092.INIT = 16'h5555;
    X_LUT4 C19092(
      .ADR0 (ADR_O[2]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12692)
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C4/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C3/C2/O ),
      .I1 (N12692),
      .O (\bridge/pci_target_unit/wishbone_master/N2985/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C4/C2 (
      .IA (ADR_O[2]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C3/C2/O ),
      .SEL (N12692),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C4/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2985/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2985/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N2986 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2985/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2985/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2985 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2985/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2985/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C5/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C7/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C6/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2987/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2987/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C7/C2 (
      .IA (ADR_O[5]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C6/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2987/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2987/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2987/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2987/G (
      .ADR0 (ADR_O[5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2987/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2987/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2987/F (
      .ADR0 (ADR_O[4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2987/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C6/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C5/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2987/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2987/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C6/C2 (
      .IA (ADR_O[4]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C5/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2987/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C6/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2987/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2987/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N2988 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2987/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2987/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2987 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2987/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2987/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C7/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C9/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C8/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2989/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2989/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C9/C2 (
      .IA (ADR_O[7]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C8/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2989/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2989/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2989/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2989/G (
      .ADR0 (ADR_O[7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2989/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2989/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2989/F (
      .ADR0 (ADR_O[6]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2989/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C8/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C7/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2989/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2989/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C8/C2 (
      .IA (ADR_O[6]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C7/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2989/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C8/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2989/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2989/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N2990 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2989/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2989/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2989 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2989/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2989/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C9/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C11/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C10/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2991/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2991/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C11/C2 (
      .IA (ADR_O[9]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C10/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2991/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2991/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2991/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2991/G (
      .ADR0 (ADR_O[9]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2991/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2991/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2991/F (
      .ADR0 (ADR_O[8]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2991/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C10/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C9/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2991/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2991/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C10/C2 (
      .IA (ADR_O[8]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C9/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2991/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C10/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2991/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2991/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N2992 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2991/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2991/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2991 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2991/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2991/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C11/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C13/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C12/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2993/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2993/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C13/C2 (
      .IA (\bridge/pciu_err_addr_out[11] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C12/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2993/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2993/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2993/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2993/G (
      .ADR0 (\bridge/pciu_err_addr_out[11] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2993/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2993/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2993/F (
      .ADR0 (ADR_O[10]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2993/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C12/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C11/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2993/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2993/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C12/C2 (
      .IA (ADR_O[10]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C11/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2993/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C12/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2993/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2993/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N2994 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2993/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2993/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2993 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2993/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2993/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C13/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C15/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C14/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2995/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2995/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C15/C2 (
      .IA (\bridge/pciu_err_addr_out[13] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C14/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2995/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2995/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2995/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2995/G (
      .ADR0 (\bridge/pciu_err_addr_out[13] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2995/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2995/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2995/F (
      .ADR0 (\bridge/pciu_err_addr_out[12] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2995/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C14/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C13/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2995/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2995/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C14/C2 (
      .IA (\bridge/pciu_err_addr_out[12] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C13/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2995/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C14/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2995/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2995/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N2996 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2995/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2995/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2995 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2995/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2995/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C15/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C17/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C16/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2997/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2997/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C17/C2 (
      .IA (\bridge/pciu_err_addr_out[15] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C16/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2997/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2997/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2997/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2997/G (
      .ADR0 (\bridge/pciu_err_addr_out[15] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2997/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2997/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2997/F (
      .ADR0 (\bridge/pciu_err_addr_out[14] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2997/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C16/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C15/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2997/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2997/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C16/C2 (
      .IA (\bridge/pciu_err_addr_out[14] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C15/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2997/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C16/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2997/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2997/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N2998 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2997/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2997/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2997 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2997/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2997/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C17/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C19/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C18/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2999/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2999/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C19/C2 (
      .IA (\bridge/pciu_err_addr_out[17] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C18/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2999/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2999/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2999/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2999/G (
      .ADR0 (\bridge/pciu_err_addr_out[17] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2999/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N2999/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N2999/F (
      .ADR0 (\bridge/pciu_err_addr_out[16] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N2999/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C18/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C17/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N2999/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N2999/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C18/C2 (
      .IA (\bridge/pciu_err_addr_out[16] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C17/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N2999/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C18/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2999/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2999/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3000 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2999/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2999/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N2999 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N2999/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N2999/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C19/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C21/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C20/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3001/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3001/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C21/C2 (
      .IA (\bridge/pciu_err_addr_out[19] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C20/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3001/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3001/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3001/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3001/G (
      .ADR0 (\bridge/pciu_err_addr_out[19] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3001/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3001/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3001/F (
      .ADR0 (\bridge/pciu_err_addr_out[18] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3001/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C20/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C19/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3001/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3001/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C20/C2 (
      .IA (\bridge/pciu_err_addr_out[18] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C19/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3001/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C20/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3001/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3001/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3002 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3001/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3001/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3001 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3001/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3001/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C21/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C23/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C22/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3003/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3003/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C23/C2 (
      .IA (\bridge/pciu_err_addr_out[21] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C22/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3003/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3003/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3003/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3003/G (
      .ADR0 (\bridge/pciu_err_addr_out[21] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3003/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3003/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3003/F (
      .ADR0 (\bridge/pciu_err_addr_out[20] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3003/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C22/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C21/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3003/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3003/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C22/C2 (
      .IA (\bridge/pciu_err_addr_out[20] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C21/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3003/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C22/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3003/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3003/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3004 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3003/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3003/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3003 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3003/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3003/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C23/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C25/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C24/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3005/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3005/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C25/C2 (
      .IA (\bridge/pciu_err_addr_out[23] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C24/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3005/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3005/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3005/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3005/G (
      .ADR0 (\bridge/pciu_err_addr_out[23] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3005/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3005/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3005/F (
      .ADR0 (\bridge/pciu_err_addr_out[22] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3005/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C24/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C23/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3005/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3005/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C24/C2 (
      .IA (\bridge/pciu_err_addr_out[22] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C23/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3005/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C24/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3005/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3005/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3006 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3005/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3005/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3005 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3005/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3005/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C25/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C27/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C26/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3007/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3007/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C27/C2 (
      .IA (\bridge/pciu_err_addr_out[25] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C26/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3007/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3007/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3007/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3007/G (
      .ADR0 (\bridge/pciu_err_addr_out[25] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3007/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3007/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3007/F (
      .ADR0 (\bridge/pciu_err_addr_out[24] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3007/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C26/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C25/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3007/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3007/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C26/C2 (
      .IA (\bridge/pciu_err_addr_out[24] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C25/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3007/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C26/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3007/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3007/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3008 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3007/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3007/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3007 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3007/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3007/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C27/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C29/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C28/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3009/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3009/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C29/C2 (
      .IA (\bridge/pciu_err_addr_out[27] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C28/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3009/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3009/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3009/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3009/G (
      .ADR0 (\bridge/pciu_err_addr_out[27] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3009/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3009/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3009/F (
      .ADR0 (\bridge/pciu_err_addr_out[26] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3009/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C28/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C27/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3009/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3009/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C28/C2 (
      .IA (\bridge/pciu_err_addr_out[26] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C27/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3009/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C28/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3009/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3009/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3010 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3009/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3009/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3009 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3009/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3009/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C29/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C31/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C30/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3011/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3011/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C31/C2 (
      .IA (\bridge/pciu_err_addr_out[29] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C30/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3011/GROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3011/CYMUXG )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3011/G .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3011/G (
      .ADR0 (\bridge/pciu_err_addr_out[29] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3011/GROM )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3011/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3011/F (
      .ADR0 (\bridge/pciu_err_addr_out[28] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3011/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C30/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C29/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3011/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3011/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C30/C2 (
      .IA (\bridge/pciu_err_addr_out[28] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C29/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3011/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C30/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3011/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3011/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3012 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3011/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3011/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3011 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3011/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3011/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C31/C2/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C33/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C32/C2/O ),
      .I1 (\bridge/pciu_err_addr_out[31]_rt ),
      .O (\bridge/pci_target_unit/wishbone_master/N3013/XORG )
    );
    defparam \bridge/pciu_err_addr_out<31>_rt .INIT = 16'hAAAA;
    X_LUT4 \bridge/pciu_err_addr_out<31>_rt (
      .ADR0 (\bridge/pciu_err_addr_out[31] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pciu_err_addr_out[31]_rt )
    );
    defparam \bridge/pci_target_unit/wishbone_master/N3013/F .INIT = 16'hAAAA;
    X_LUT4 \bridge/pci_target_unit/wishbone_master/N3013/F (
      .ADR0 (\bridge/pciu_err_addr_out[30] ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/N3013/FROM )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3409/C32/C1 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3409/C31/C2/O ),
      .I1 (\bridge/pci_target_unit/wishbone_master/N3013/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/N3013/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3409/C32/C2 (
      .IA (\bridge/pciu_err_addr_out[30] ),
      .IB (\bridge/pci_target_unit/wishbone_master/C3409/C31/C2/O ),
      .SEL (\bridge/pci_target_unit/wishbone_master/N3013/FROM ),
      .O (\bridge/pci_target_unit/wishbone_master/C3409/C32/C2/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3013/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3013/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3014 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3013/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3013/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3013 )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3411/C4/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3411/C3/C1/O ),
      .I1 (N12696),
      .O (\bridge/pci_target_unit/wishbone_master/N3110/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3411/C4/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/cache_line [1]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3411/C3/C1/O ),
      .SEL (N12696),
      .O (\bridge/pci_target_unit/wishbone_master/N3110/CYMUXG )
    );
    defparam C19082.INIT = 16'h5555;
    X_LUT4 C19082(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [1]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12696)
    );
    defparam C19083.INIT = 16'h5555;
    X_LUT4 C19083(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [0]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12694)
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3411/C3/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/N3110/LOGIC_ZERO ),
      .I1 (N12694),
      .O (\bridge/pci_target_unit/wishbone_master/N3110/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3411/C3/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/cache_line [0]),
      .IB (\bridge/pci_target_unit/wishbone_master/N3110/LOGIC_ZERO ),
      .SEL (N12694),
      .O (\bridge/pci_target_unit/wishbone_master/C3411/C3/C1/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3110/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3110/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3111 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3110/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3110/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3110 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3110/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3110/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3411/C4/C1/O )
    );
    X_ZERO \bridge/pci_target_unit/wishbone_master/N3110/LOGIC_ZERO_301 (
      .O (\bridge/pci_target_unit/wishbone_master/N3110/LOGIC_ZERO )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3411/C6/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3411/C5/C1/O ),
      .I1 (N12700),
      .O (\bridge/pci_target_unit/wishbone_master/N3112/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3411/C6/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/cache_line [3]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3411/C5/C1/O ),
      .SEL (N12700),
      .O (\bridge/pci_target_unit/wishbone_master/N3112/CYMUXG )
    );
    defparam C19080.INIT = 16'h5555;
    X_LUT4 C19080(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12700)
    );
    defparam C19081.INIT = 16'h5555;
    X_LUT4 C19081(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [2]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12698)
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3411/C5/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3411/C4/C1/O ),
      .I1 (N12698),
      .O (\bridge/pci_target_unit/wishbone_master/N3112/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3411/C5/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/cache_line [2]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3411/C4/C1/O ),
      .SEL (N12698),
      .O (\bridge/pci_target_unit/wishbone_master/C3411/C5/C1/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3112/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3112/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3113 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3112/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3112/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3112 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3112/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3112/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3411/C6/C1/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3411/C8/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3411/C7/C1/O ),
      .I1 (N12704),
      .O (\bridge/pci_target_unit/wishbone_master/N3114/XORG )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3411/C8/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/cache_line [5]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3411/C7/C1/O ),
      .SEL (N12704),
      .O (\bridge/pci_target_unit/wishbone_master/N3114/CYMUXG )
    );
    defparam C19078.INIT = 16'h5555;
    X_LUT4 C19078(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12704)
    );
    defparam C19079.INIT = 16'h5555;
    X_LUT4 C19079(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12702)
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3411/C7/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3411/C6/C1/O ),
      .I1 (N12702),
      .O (\bridge/pci_target_unit/wishbone_master/N3114/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3411/C7/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/cache_line [4]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3411/C6/C1/O ),
      .SEL (N12702),
      .O (\bridge/pci_target_unit/wishbone_master/C3411/C7/C1/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3114/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3114/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3115 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3114/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3114/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3114 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3114/COUTUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3114/CYMUXG ),
      .O (\bridge/pci_target_unit/wishbone_master/C3411/C8/C1/O )
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3411/C10/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3411/C9/C1/O ),
      .I1 (N12708),
      .O (\bridge/pci_target_unit/wishbone_master/N3116/XORG )
    );
    defparam C19076.INIT = 16'h5555;
    X_LUT4 C19076(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12708)
    );
    defparam C19077.INIT = 16'h5555;
    X_LUT4 C19077(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/cache_line [6]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12706)
    );
    X_XOR2 \bridge/pci_target_unit/wishbone_master/C3411/C9/C0 (
      .I0 (\bridge/pci_target_unit/wishbone_master/C3411/C8/C1/O ),
      .I1 (N12706),
      .O (\bridge/pci_target_unit/wishbone_master/N3116/XORF )
    );
    X_MUX2 \bridge/pci_target_unit/wishbone_master/C3411/C9/C1 (
      .IA (\bridge/pci_target_unit/wishbone_master/cache_line [6]),
      .IB (\bridge/pci_target_unit/wishbone_master/C3411/C8/C1/O ),
      .SEL (N12706),
      .O (\bridge/pci_target_unit/wishbone_master/C3411/C9/C1/O )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3116/YUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3116/XORG ),
      .O (\bridge/pci_target_unit/wishbone_master/N3117 )
    );
    X_BUF \bridge/pci_target_unit/wishbone_master/N3116/XUSED (
      .I (\bridge/pci_target_unit/wishbone_master/N3116/XORF ),
      .O (\bridge/pci_target_unit/wishbone_master/N3116 )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C4/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C3/C1/O ),
      .I1 (N12657),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C4/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [1]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C3/C1/O ),
      .SEL (N12657),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/CYMUXG )
    );
    defparam C19108.INIT = 16'h5555;
    X_LUT4 C19108(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [1]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12657)
    );
    defparam C19109.INIT = 16'h5555;
    X_LUT4 C19109(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [0]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12655)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C3/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/LOGIC_ZERO ),
      .I1 (N12655),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C3/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [0]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/LOGIC_ZERO ),
      .SEL (N12655),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C3/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2618/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2619 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2618/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2618/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C4/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_sm/N2618/LOGIC_ZERO_302 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2618/LOGIC_ZERO )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C6/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C5/C1/O ),
      .I1 (N12661),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2620/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C6/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [3]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C5/C1/O ),
      .SEL (N12661),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2620/CYMUXG )
    );
    defparam C19106.INIT = 16'h5555;
    X_LUT4 C19106(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12661)
    );
    defparam C19107.INIT = 16'h5555;
    X_LUT4 C19107(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [2]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12659)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C5/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C4/C1/O ),
      .I1 (N12659),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2620/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C5/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [2]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C4/C1/O ),
      .SEL (N12659),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C5/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2620/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2620/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2621 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2620/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2620/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2620 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2620/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2620/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C6/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C8/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C7/C1/O ),
      .I1 (N12665),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2622/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C8/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [5]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C7/C1/O ),
      .SEL (N12665),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2622/CYMUXG )
    );
    defparam C19104.INIT = 16'h5555;
    X_LUT4 C19104(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12665)
    );
    defparam C19105.INIT = 16'h5555;
    X_LUT4 C19105(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12663)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C7/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C6/C1/O ),
      .I1 (N12663),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2622/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C7/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [4]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C6/C1/O ),
      .SEL (N12663),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C7/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2622/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2622/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2623 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2622/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2622/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2622 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2622/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2622/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C8/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C10/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C9/C1/O ),
      .I1 (N12669),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2624/XORG )
    );
    defparam C19102.INIT = 16'h5555;
    X_LUT4 C19102(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12669)
    );
    defparam C19103.INIT = 16'h5555;
    X_LUT4 C19103(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [6]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12667)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C9/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C8/C1/O ),
      .I1 (N12667),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2624/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C9/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_sm/latency_timer [6]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C8/C1/O ),
      .SEL (N12667),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/C2703/C9/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2624/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2624/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2625 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_sm/N2624/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_sm/N2624/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_sm/N2624 )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C4/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C3/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N140/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N140/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C4/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C3/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N140/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N140/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N140/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N140/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [1]),
      .O (\bridge/wishbone_slave_unit/del_sync/N140/GROM )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N140/F .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N140/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [0]),
      .O (\bridge/wishbone_slave_unit/del_sync/N140/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C3/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ONE ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N140/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N140/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C3/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ONE ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N140/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C3/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ZERO_303 (
      .O (\bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N140/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N140/XORG ),
      .O (\bridge/wishbone_slave_unit/del_sync/N141 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N140/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N140/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N140 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N140/COUTUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N140/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C4/C1/O )
    );
    X_ONE \bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ONE_304 (
      .O (\bridge/wishbone_slave_unit/del_sync/N140/LOGIC_ONE )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C6/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C5/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N142/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N142/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C6/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N142/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C5/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N142/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N142/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N142/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N142/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [3]),
      .O (\bridge/wishbone_slave_unit/del_sync/N142/GROM )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N142/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N142/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [2]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/N142/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C5/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C4/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N142/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N142/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C5/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N142/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C4/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N142/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C5/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/del_sync/N142/LOGIC_ZERO_305 (
      .O (\bridge/wishbone_slave_unit/del_sync/N142/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N142/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N142/XORG ),
      .O (\bridge/wishbone_slave_unit/del_sync/N143 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N142/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N142/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N142 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N142/COUTUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N142/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C6/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C8/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C7/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N144/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N144/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C8/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N144/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C7/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N144/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N144/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N144/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N144/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [5]),
      .O (\bridge/wishbone_slave_unit/del_sync/N144/GROM )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N144/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N144/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [4]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/N144/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C7/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C6/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N144/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N144/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C7/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N144/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C6/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N144/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C7/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/del_sync/N144/LOGIC_ZERO_306 (
      .O (\bridge/wishbone_slave_unit/del_sync/N144/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N144/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N144/XORG ),
      .O (\bridge/wishbone_slave_unit/del_sync/N145 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N144/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N144/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N144 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N144/COUTUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N144/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C8/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C10/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C9/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N146/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N146/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C10/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N146/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C9/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N146/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N146/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N146/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N146/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [7]),
      .O (\bridge/wishbone_slave_unit/del_sync/N146/GROM )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N146/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N146/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [6]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/N146/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C9/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C8/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N146/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N146/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C9/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N146/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C8/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N146/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C9/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/del_sync/N146/LOGIC_ZERO_307 (
      .O (\bridge/wishbone_slave_unit/del_sync/N146/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N146/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N146/XORG ),
      .O (\bridge/wishbone_slave_unit/del_sync/N147 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N146/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N146/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N146 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N146/COUTUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N146/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C10/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C12/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C11/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N148/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N148/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C12/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N148/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C11/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N148/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N148/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N148/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N148/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [9]),
      .O (\bridge/wishbone_slave_unit/del_sync/N148/GROM )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N148/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N148/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [8]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/N148/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C11/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C10/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N148/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N148/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C11/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N148/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C10/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N148/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C11/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/del_sync/N148/LOGIC_ZERO_308 (
      .O (\bridge/wishbone_slave_unit/del_sync/N148/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N148/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N148/XORG ),
      .O (\bridge/wishbone_slave_unit/del_sync/N149 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N148/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N148/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N148 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N148/COUTUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N148/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C12/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C14/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C13/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N150/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N150/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C14/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N150/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C13/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N150/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N150/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N150/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N150/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [11]),
      .O (\bridge/wishbone_slave_unit/del_sync/N150/GROM )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N150/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N150/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [10]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/N150/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C13/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C12/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N150/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N150/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C13/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N150/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C12/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N150/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C13/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/del_sync/N150/LOGIC_ZERO_309 (
      .O (\bridge/wishbone_slave_unit/del_sync/N150/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N150/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N150/XORG ),
      .O (\bridge/wishbone_slave_unit/del_sync/N151 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N150/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N150/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N150 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N150/COUTUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N150/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C14/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C16/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C15/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N152/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N152/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C16/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N152/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C15/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N152/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N152/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N152/G .INIT = 16'hCCCC;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N152/G (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [13]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/N152/GROM )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N152/F .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N152/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [12]),
      .O (\bridge/wishbone_slave_unit/del_sync/N152/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C15/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C14/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N152/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N152/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C15/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N152/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C14/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N152/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C15/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/del_sync/N152/LOGIC_ZERO_310 (
      .O (\bridge/wishbone_slave_unit/del_sync/N152/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N152/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N152/XORG ),
      .O (\bridge/wishbone_slave_unit/del_sync/N153 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N152/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N152/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N152 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N152/COUTUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N152/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C16/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C18/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C17/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N154/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N154/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C18/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N154/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C17/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N154/GROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N154/CYMUXG )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N154/G .INIT = 16'hFF00;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N154/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [15]),
      .O (\bridge/wishbone_slave_unit/del_sync/N154/GROM )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/N154/F .INIT = 16'hF0F0;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/N154/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [14]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/N154/FROM )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C17/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C16/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/N154/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/N154/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/del_sync/C24/C17/C1 (
      .IA (\bridge/wishbone_slave_unit/del_sync/N154/LOGIC_ZERO ),
      .IB (\bridge/wishbone_slave_unit/del_sync/C24/C16/C1/O ),
      .SEL (\bridge/wishbone_slave_unit/del_sync/N154/FROM ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C17/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/del_sync/N154/LOGIC_ZERO_311 (
      .O (\bridge/wishbone_slave_unit/del_sync/N154/LOGIC_ZERO )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N154/YUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N154/XORG ),
      .O (\bridge/wishbone_slave_unit/del_sync/N155 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N154/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N154/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N154 )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N154/COUTUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N154/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/del_sync/C24/C18/C1/O )
    );
    defparam \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<16>_rt .INIT = 16'hCCCC;
    X_LUT4 \bridge/wishbone_slave_unit/del_sync/comp_cycle_count<16>_rt (
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count [16]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[16]_rt )
    );
    X_XOR2 \bridge/wishbone_slave_unit/del_sync/C24/C19/C0 (
      .I0 (\bridge/wishbone_slave_unit/del_sync/C24/C18/C1/O ),
      .I1 (\bridge/wishbone_slave_unit/del_sync/comp_cycle_count[16]_rt ),
      .O (\bridge/wishbone_slave_unit/del_sync/N156/XORF )
    );
    X_BUF \bridge/wishbone_slave_unit/del_sync/N156/XUSED (
      .I (\bridge/wishbone_slave_unit/del_sync/N156/XORF ),
      .O (\bridge/wishbone_slave_unit/del_sync/N156 )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C4/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C3/C1/O ),
      .I1 (\CRT/ssvga_crtc/N400/GROM ),
      .O (\CRT/ssvga_crtc/N400/XORG )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C4/C1 (
      .IA (\CRT/ssvga_crtc/N400/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C530/C3/C1/O ),
      .SEL (\CRT/ssvga_crtc/N400/GROM ),
      .O (\CRT/ssvga_crtc/N400/CYMUXG )
    );
    defparam \CRT/ssvga_crtc/N400/G .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_crtc/N400/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/hcntr [1]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N400/GROM )
    );
    defparam \CRT/ssvga_crtc/N400/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_crtc/N400/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/hcntr [0]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N400/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C3/C0 (
      .I0 (\CRT/ssvga_crtc/N400/LOGIC_ONE ),
      .I1 (\CRT/ssvga_crtc/N400/FROM ),
      .O (\CRT/ssvga_crtc/N400/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C3/C1 (
      .IA (\CRT/ssvga_crtc/N400/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/N400/LOGIC_ONE ),
      .SEL (\CRT/ssvga_crtc/N400/FROM ),
      .O (\CRT/ssvga_crtc/C530/C3/C1/O )
    );
    X_ZERO \CRT/ssvga_crtc/N400/LOGIC_ZERO_312 (
      .O (\CRT/ssvga_crtc/N400/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_crtc/N400/YUSED (
      .I (\CRT/ssvga_crtc/N400/XORG ),
      .O (\CRT/ssvga_crtc/N401 )
    );
    X_BUF \CRT/ssvga_crtc/N400/XUSED (
      .I (\CRT/ssvga_crtc/N400/XORF ),
      .O (\CRT/ssvga_crtc/N400 )
    );
    X_BUF \CRT/ssvga_crtc/N400/COUTUSED (
      .I (\CRT/ssvga_crtc/N400/CYMUXG ),
      .O (\CRT/ssvga_crtc/C530/C4/C1/O )
    );
    X_ONE \CRT/ssvga_crtc/N400/LOGIC_ONE_313 (
      .O (\CRT/ssvga_crtc/N400/LOGIC_ONE )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C6/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C5/C1/O ),
      .I1 (\CRT/ssvga_crtc/N402/GROM ),
      .O (\CRT/ssvga_crtc/N402/XORG )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C6/C1 (
      .IA (\CRT/ssvga_crtc/N402/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C530/C5/C1/O ),
      .SEL (\CRT/ssvga_crtc/N402/GROM ),
      .O (\CRT/ssvga_crtc/N402/CYMUXG )
    );
    defparam \CRT/ssvga_crtc/N402/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_crtc/N402/G (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/hcntr [3]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N402/GROM )
    );
    defparam \CRT/ssvga_crtc/N402/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_crtc/N402/F (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/hcntr [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N402/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C5/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C4/C1/O ),
      .I1 (\CRT/ssvga_crtc/N402/FROM ),
      .O (\CRT/ssvga_crtc/N402/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C5/C1 (
      .IA (\CRT/ssvga_crtc/N402/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C530/C4/C1/O ),
      .SEL (\CRT/ssvga_crtc/N402/FROM ),
      .O (\CRT/ssvga_crtc/C530/C5/C1/O )
    );
    X_ZERO \CRT/ssvga_crtc/N402/LOGIC_ZERO_314 (
      .O (\CRT/ssvga_crtc/N402/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_crtc/N402/YUSED (
      .I (\CRT/ssvga_crtc/N402/XORG ),
      .O (\CRT/ssvga_crtc/N403 )
    );
    X_BUF \CRT/ssvga_crtc/N402/XUSED (
      .I (\CRT/ssvga_crtc/N402/XORF ),
      .O (\CRT/ssvga_crtc/N402 )
    );
    X_BUF \CRT/ssvga_crtc/N402/COUTUSED (
      .I (\CRT/ssvga_crtc/N402/CYMUXG ),
      .O (\CRT/ssvga_crtc/C530/C6/C1/O )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C8/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C7/C1/O ),
      .I1 (\CRT/ssvga_crtc/N404/GROM ),
      .O (\CRT/ssvga_crtc/N404/XORG )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C8/C1 (
      .IA (\CRT/ssvga_crtc/N404/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C530/C7/C1/O ),
      .SEL (\CRT/ssvga_crtc/N404/GROM ),
      .O (\CRT/ssvga_crtc/N404/CYMUXG )
    );
    defparam \CRT/ssvga_crtc/N404/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_crtc/N404/G (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/hcntr [5]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N404/GROM )
    );
    defparam \CRT/ssvga_crtc/N404/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_crtc/N404/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/hcntr [4]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N404/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C7/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C6/C1/O ),
      .I1 (\CRT/ssvga_crtc/N404/FROM ),
      .O (\CRT/ssvga_crtc/N404/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C7/C1 (
      .IA (\CRT/ssvga_crtc/N404/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C530/C6/C1/O ),
      .SEL (\CRT/ssvga_crtc/N404/FROM ),
      .O (\CRT/ssvga_crtc/C530/C7/C1/O )
    );
    X_ZERO \CRT/ssvga_crtc/N404/LOGIC_ZERO_315 (
      .O (\CRT/ssvga_crtc/N404/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_crtc/N404/YUSED (
      .I (\CRT/ssvga_crtc/N404/XORG ),
      .O (\CRT/ssvga_crtc/N405 )
    );
    X_BUF \CRT/ssvga_crtc/N404/XUSED (
      .I (\CRT/ssvga_crtc/N404/XORF ),
      .O (\CRT/ssvga_crtc/N404 )
    );
    X_BUF \CRT/ssvga_crtc/N404/COUTUSED (
      .I (\CRT/ssvga_crtc/N404/CYMUXG ),
      .O (\CRT/ssvga_crtc/C530/C8/C1/O )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C10/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C9/C1/O ),
      .I1 (\CRT/ssvga_crtc/N406/GROM ),
      .O (\CRT/ssvga_crtc/N406/XORG )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C10/C1 (
      .IA (\CRT/ssvga_crtc/N406/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C530/C9/C1/O ),
      .SEL (\CRT/ssvga_crtc/N406/GROM ),
      .O (\CRT/ssvga_crtc/N406/CYMUXG )
    );
    defparam \CRT/ssvga_crtc/N406/G .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_crtc/N406/G (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/hcntr [7]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N406/GROM )
    );
    defparam \CRT/ssvga_crtc/N406/F .INIT = 16'hF0F0;
    X_LUT4 \CRT/ssvga_crtc/N406/F (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\CRT/ssvga_crtc/hcntr [6]),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N406/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C9/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C8/C1/O ),
      .I1 (\CRT/ssvga_crtc/N406/FROM ),
      .O (\CRT/ssvga_crtc/N406/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C9/C1 (
      .IA (\CRT/ssvga_crtc/N406/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C530/C8/C1/O ),
      .SEL (\CRT/ssvga_crtc/N406/FROM ),
      .O (\CRT/ssvga_crtc/C530/C9/C1/O )
    );
    X_ZERO \CRT/ssvga_crtc/N406/LOGIC_ZERO_316 (
      .O (\CRT/ssvga_crtc/N406/LOGIC_ZERO )
    );
    X_BUF \CRT/ssvga_crtc/N406/YUSED (
      .I (\CRT/ssvga_crtc/N406/XORG ),
      .O (\CRT/ssvga_crtc/N407 )
    );
    X_BUF \CRT/ssvga_crtc/N406/XUSED (
      .I (\CRT/ssvga_crtc/N406/XORF ),
      .O (\CRT/ssvga_crtc/N406 )
    );
    X_BUF \CRT/ssvga_crtc/N406/COUTUSED (
      .I (\CRT/ssvga_crtc/N406/CYMUXG ),
      .O (\CRT/ssvga_crtc/C530/C10/C1/O )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C12/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C11/C1/O ),
      .I1 (\CRT/ssvga_crtc/hcntr[9]_rt ),
      .O (\CRT/ssvga_crtc/N408/XORG )
    );
    defparam \CRT/ssvga_crtc/hcntr<9>_rt .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_crtc/hcntr<9>_rt (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/hcntr [9]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/hcntr[9]_rt )
    );
    defparam \CRT/ssvga_crtc/N408/F .INIT = 16'hCCCC;
    X_LUT4 \CRT/ssvga_crtc/N408/F (
      .ADR0 (VCC),
      .ADR1 (\CRT/ssvga_crtc/hcntr [8]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\CRT/ssvga_crtc/N408/FROM )
    );
    X_XOR2 \CRT/ssvga_crtc/C530/C11/C0 (
      .I0 (\CRT/ssvga_crtc/C530/C10/C1/O ),
      .I1 (\CRT/ssvga_crtc/N408/FROM ),
      .O (\CRT/ssvga_crtc/N408/XORF )
    );
    X_MUX2 \CRT/ssvga_crtc/C530/C11/C1 (
      .IA (\CRT/ssvga_crtc/N408/LOGIC_ZERO ),
      .IB (\CRT/ssvga_crtc/C530/C10/C1/O ),
      .SEL (\CRT/ssvga_crtc/N408/FROM ),
      .O (\CRT/ssvga_crtc/C530/C11/C1/O )
    );
    X_BUF \CRT/ssvga_crtc/N408/YUSED (
      .I (\CRT/ssvga_crtc/N408/XORG ),
      .O (\CRT/ssvga_crtc/N409 )
    );
    X_BUF \CRT/ssvga_crtc/N408/XUSED (
      .I (\CRT/ssvga_crtc/N408/XORF ),
      .O (\CRT/ssvga_crtc/N408 )
    );
    X_ZERO \CRT/ssvga_crtc/N408/LOGIC_ZERO_317 (
      .O (\CRT/ssvga_crtc/N408/LOGIC_ZERO )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C4/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C3/C1/O ),
      .I1 (N12675),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C4/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [1]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C3/C1/O ),
      .SEL (N12675),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/CYMUXG )
    );
    defparam C19100.INIT = 16'h5555;
    X_LUT4 C19100(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [1]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12675)
    );
    defparam C19101.INIT = 16'h5555;
    X_LUT4 C19101(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [0]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12673)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C3/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/LOGIC_ZERO ),
      .I1 (N12673),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C3/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [0]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/LOGIC_ZERO ),
      .SEL (N12673),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C3/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3190/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3191 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3190/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3190 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3190/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C4/C1/O )
    );
    X_ZERO \bridge/wishbone_slave_unit/pci_initiator_if/N3190/LOGIC_ZERO_318 (
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3190/LOGIC_ZERO )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C6/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C5/C1/O ),
      .I1 (N12679),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3192/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C6/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [3]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C5/C1/O ),
      .SEL (N12679),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3192/CYMUXG )
    );
    defparam C19098.INIT = 16'h5555;
    X_LUT4 C19098(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [3]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12679)
    );
    defparam C19099.INIT = 16'h5555;
    X_LUT4 C19099(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [2]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12677)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C5/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C4/C1/O ),
      .I1 (N12677),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3192/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C5/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [2]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C4/C1/O ),
      .SEL (N12677),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C5/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3192/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3192/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3193 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3192/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3192/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3192 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3192/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3192/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C6/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C8/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C7/C1/O ),
      .I1 (N12683),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3194/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C8/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [5]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C7/C1/O ),
      .SEL (N12683),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3194/CYMUXG )
    );
    defparam C19096.INIT = 16'h5555;
    X_LUT4 C19096(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [5]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12683)
    );
    defparam C19097.INIT = 16'h5555;
    X_LUT4 C19097(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [4]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12681)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C7/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C6/C1/O ),
      .I1 (N12681),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3194/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C7/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [4]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C6/C1/O ),
      .SEL (N12681),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C7/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3194/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3194/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3195 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3194/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3194/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3194 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3194/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3194/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C8/C1/O )
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C10/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C9/C1/O ),
      .I1 (N12687),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3196/XORG )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C10/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [7]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C9/C1/O ),
      .SEL (N12687),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3196/CYMUXG )
    );
    defparam C19094.INIT = 16'h5555;
    X_LUT4 C19094(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [7]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12687)
    );
    defparam C19095.INIT = 16'h5555;
    X_LUT4 C19095(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [6]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12685)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C9/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C8/C1/O ),
      .I1 (N12685),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3196/XORF )
    );
    X_MUX2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C9/C1 (
      .IA (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [6]),
      .IB (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C8/C1/O ),
      .SEL (N12685),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C9/C1/O )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3196/YUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3196/XORG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3197 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3196/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3196/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3196 )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3196/COUTUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3196/CYMUXG ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C10/C1/O )
    );
    defparam C19093.INIT = 16'h5555;
    X_LUT4 C19093(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/read_count [8]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (N12689)
    );
    X_XOR2 \bridge/wishbone_slave_unit/pci_initiator_if/C3273/C11/C0 (
      .I0 (\bridge/wishbone_slave_unit/pci_initiator_if/C3273/C10/C1/O ),
      .I1 (N12689),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3198/XORF )
    );
    X_BUF \bridge/wishbone_slave_unit/pci_initiator_if/N3198/XUSED (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/N3198/XORF ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/N3198 )
    );
    defparam C18412.INIT = 16'hFE02;
    X_LUT4 C18412(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [24]),
      .ADR1 (\bridge/in_reg_trdy_out ),
      .ADR2 (\bridge/in_reg_devsel_out ),
      .ADR3 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [24]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/GROM )
    );
    defparam C18395.INIT = 16'hCCCA;
    X_LUT4 C18395(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [25]),
      .ADR1 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [25]),
      .ADR2 (\bridge/in_reg_trdy_out ),
      .ADR3 (\bridge/in_reg_devsel_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<25>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<25>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [24])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<25>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [25])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<24> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [24])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<25> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [25])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[25]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18538.INIT = 16'hAFA0;
    X_LUT4 C18538(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [16]),
      .ADR1 (VCC),
      .ADR2 (syn18908),
      .ADR3 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [16]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/GROM )
    );
    defparam C18522.INIT = 16'hAACC;
    X_LUT4 C18522(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [17]),
      .ADR1 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [17]),
      .ADR2 (VCC),
      .ADR3 (syn18908),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<17>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<17>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [16])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<17>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [17])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<16> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [16])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<17> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [17])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[17]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18036.INIT = 16'h2222;
    X_LUT4 C18036(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [30]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N12 )
    );
    defparam C18035.INIT = 16'h5500;
    X_LUT4 C18035(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [31]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N6 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<31>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<30> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [30])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<31>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<31> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [31])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<31>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[31]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18044.INIT = 16'h5050;
    X_LUT4 C18044(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [22]),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N60 )
    );
    defparam C18043.INIT = 16'h5500;
    X_LUT4 C18043(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [23]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N54 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<23>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<22> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N60 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [22])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<23>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<23> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N54 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [23])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<23>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[23]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18052.INIT = 16'h2222;
    X_LUT4 C18052(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [14]),
      .ADR1 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N108 )
    );
    defparam C18051.INIT = 16'h5500;
    X_LUT4 C18051(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [15]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N102 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<15>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<14> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N108 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [14])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<15>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<15> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N102 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [15])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<15>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[15]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17823.INIT = 16'hFCB8;
    X_LUT4 C17823(
      .ADR0 (\bridge/conf_cache_line_size_out [0]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/N3110 ),
      .ADR3 (syn23022),
      .O (\bridge/pci_target_unit/wishbone_master/C3414/N6 )
    );
    defparam C17821.INIT = 16'hBB88;
    X_LUT4 C17821(
      .ADR0 (\bridge/conf_cache_line_size_out [1]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/N3111 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3414/N12 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/cache_line<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line[1]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/cache_line_reg<0> (
      .I (\bridge/pci_target_unit/wishbone_master/C3414/N6 ),
      .CLK (CLK_BUFGPed),
      .CE (N12510),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/cache_line[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line [0])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/cache_line<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/cache_line[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/cache_line[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/cache_line_reg<1> (
      .I (\bridge/pci_target_unit/wishbone_master/C3414/N12 ),
      .CLK (CLK_BUFGPed),
      .CE (N12510),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/cache_line[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line [1])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/cache_line<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/cache_line[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/cache_line[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18378.INIT = 16'hF0E4;
    X_LUT4 C18378(
      .ADR0 (\bridge/in_reg_devsel_out ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [26]),
      .ADR2 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [26]),
      .ADR3 (\bridge/in_reg_trdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/GROM )
    );
    defparam C18361.INIT = 16'hF0E2;
    X_LUT4 C18361(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [27]),
      .ADR1 (\bridge/in_reg_devsel_out ),
      .ADR2 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [27]),
      .ADR3 (\bridge/in_reg_trdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<27>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<27>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [26])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<27>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [27])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<26> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [26])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<27> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [27])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[27]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18506.INIT = 16'hFE10;
    X_LUT4 C18506(
      .ADR0 (\bridge/in_reg_devsel_out ),
      .ADR1 (\bridge/in_reg_trdy_out ),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [18]),
      .ADR3 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [18]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/GROM )
    );
    defparam C18491.INIT = 16'hF0E2;
    X_LUT4 C18491(
      .ADR0 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [19]),
      .ADR1 (\bridge/in_reg_devsel_out ),
      .ADR2 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [19]),
      .ADR3 (\bridge/in_reg_trdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<19>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<19>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [18])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<19>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [19])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<18> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [18])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<19> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [19])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[19]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18042.INIT = 16'h4444;
    X_LUT4 C18042(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [24]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N48 )
    );
    defparam C18041.INIT = 16'h5500;
    X_LUT4 C18041(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [25]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N42 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<25>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<24> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N48 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [24])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<25>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<25> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N42 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [25])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<25>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[25]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18050.INIT = 16'h0F00;
    X_LUT4 C18050(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [16]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N96 )
    );
    defparam C18049.INIT = 16'h0C0C;
    X_LUT4 C18049(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [17]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N90 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<17>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<16> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N96 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [16])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<17>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<17> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N90 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [17])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<17>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[17]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17820.INIT = 16'hCACA;
    X_LUT4 C17820(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3112 ),
      .ADR1 (\bridge/conf_cache_line_size_out [2]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/C3414/N18 )
    );
    defparam C17819.INIT = 16'hACAC;
    X_LUT4 C17819(
      .ADR0 (\bridge/conf_cache_line_size_out [3]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3113 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/C3414/N24 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/cache_line<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line[3]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/cache_line_reg<2> (
      .I (\bridge/pci_target_unit/wishbone_master/C3414/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (N12510),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/cache_line[3]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line [2])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/cache_line<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/cache_line[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/cache_line[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/cache_line_reg<3> (
      .I (\bridge/pci_target_unit/wishbone_master/C3414/N24 ),
      .CLK (CLK_BUFGPed),
      .CE (N12510),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/cache_line[3]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line [3])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/cache_line<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/cache_line[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/cache_line[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18342.INIT = 16'hABA8;
    X_LUT4 C18342(
      .ADR0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [28]),
      .ADR1 (\bridge/in_reg_trdy_out ),
      .ADR2 (\bridge/in_reg_devsel_out ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [28]),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/GROM )
    );
    defparam C18324.INIT = 16'hCCD8;
    X_LUT4 C18324(
      .ADR0 (\bridge/in_reg_devsel_out ),
      .ADR1 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [29]),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [29]),
      .ADR3 (\bridge/in_reg_trdy_out ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/FROM )
    );
    X_INV \bridge/wishbone_slave_unit/pcim_if_data_out<29>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<29>/YUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/GROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [28])
    );
    X_BUF \bridge/wishbone_slave_unit/pcim_if_data_out<29>/XUSED (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/FROM ),
      .O (\bridge/wishbone_slave_unit/pcim_if_next_data_out [29])
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<28> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [28])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/pci_initiator_if/data_out_reg<29> (
      .I (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/FROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/data_be_load ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out [29])
    );
    X_OR2 \bridge/wishbone_slave_unit/pcim_if_data_out<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/SRNOT ),
      .I1 (GSR),
      .O (\bridge/wishbone_slave_unit/pcim_if_data_out[29]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17659.INIT = 16'h55AA;
    X_LUT4 C17659(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [1]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_waddr [0]),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[1]/GROM )
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_waddr<1>/YUSED (
      .I (\bridge/pci_target_unit/fifos/pcir_waddr[1]/GROM ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next [0])
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next_reg<0> (
      .I (\bridge/pci_target_unit/fifos/pcir_waddr[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_waddr[1]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [0])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_waddr<1>/FFY/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[1]/FFY/RST )
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_waddr<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_waddr[1]/FFY/RST ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[1]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/waddr_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST (\bridge/pci_target_unit/fifos/pcir_waddr[1]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr [1])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_waddr<1>/FFX/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[1]/FFX/RST )
    );
    X_OR2 \bridge/pci_target_unit/fifos/pcir_waddr<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_waddr[1]/FFX/RST ),
      .I1 (GSR),
      .O (\bridge/pci_target_unit/fifos/pcir_waddr[1]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18040.INIT = 16'h00F0;
    X_LUT4 C18040(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [26]),
      .ADR3 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N36 )
    );
    defparam C18039.INIT = 16'h5500;
    X_LUT4 C18039(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [27]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N30 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<27>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<26> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [26])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<27>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<27> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [27])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<27>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[27]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18048.INIT = 16'h4444;
    X_LUT4 C18048(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [18]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N84 )
    );
    defparam C18047.INIT = 16'h5500;
    X_LUT4 C18047(
      .ADR0 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [19]),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N78 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<19>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<18> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N84 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [18])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<19>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<19> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N78 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [19])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<19>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[19]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17684.INIT = 16'h3C3C;
    X_LUT4 C17684(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_waddr [1]),
      .ADR2 (\bridge/pci_target_unit/fifos/pcir_waddr [2]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next [1])
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next_reg<1> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [1])
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_clear ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[1]/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C17818.INIT = 16'hCACA;
    X_LUT4 C17818(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3114 ),
      .ADR1 (\bridge/conf_cache_line_size_out [4]),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/C3414/N30 )
    );
    defparam C17817.INIT = 16'hE4E4;
    X_LUT4 C17817(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3115 ),
      .ADR2 (\bridge/conf_cache_line_size_out [5]),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/C3414/N36 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/cache_line<5>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line[5]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/cache_line_reg<4> (
      .I (\bridge/pci_target_unit/wishbone_master/C3414/N30 ),
      .CLK (CLK_BUFGPed),
      .CE (N12510),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/cache_line[5]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line [4])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/cache_line<5>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/cache_line[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/cache_line[5]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/cache_line_reg<5> (
      .I (\bridge/pci_target_unit/wishbone_master/C3414/N36 ),
      .CLK (CLK_BUFGPed),
      .CE (N12510),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/cache_line[5]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line [5])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/cache_line<5>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/cache_line[5]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/cache_line[5]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17663.INIT = 16'h55AA;
    X_LUT4 C17663(
      .ADR0 (\bridge/pci_target_unit/fifos/pcir_waddr [2]),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_waddr [3]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next [2])
    );
    defparam C17680.INIT = 16'h33CC;
    X_LUT4 C17680(
      .ADR0 (VCC),
      .ADR1 (\bridge/pci_target_unit/fifos/pcir_waddr [4]),
      .ADR2 (VCC),
      .ADR3 (\bridge/pci_target_unit/fifos/pcir_waddr [3]),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next [3])
    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next_reg<2> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [2])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next<3>/FFY/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFY/RST )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFY/RST ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next_reg<3> (
      .I (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/calc_wgrey_next [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next [3])
    );
    X_BUF \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next<3>/FFX/RSTOR (
      .I (\bridge/pci_target_unit/fifos/pcir_clear ),
      .O (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFX/RST )
    );
    X_OR2
     \bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFX/RST ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/fifos/pcir_fifo_ctrl/wgrey_next[3]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18038.INIT = 16'h0C0C;
    X_LUT4 C18038(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [28]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N24 )
    );
    defparam C18037.INIT = 16'h0C0C;
    X_LUT4 C18037(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [29]),
      .ADR2 (\bridge/wishbone_slave_unit/pci_initiator_if/data_source ),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N18 )
    );
    X_INV
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<29>/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/SRNOT )
    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<28> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N24 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [28])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<29>/FFY/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data_reg<29> (
      .I (\bridge/wishbone_slave_unit/pci_initiator_if/C13/N18 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_enable ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data [29])
    );
    X_OR2
     \bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data<29>/FFX/ASYNC_FF_GSR_OR (
      .I0 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/pci_initiator_if/intermediate_data[29]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C18141.INIT = 16'hCC00;
    X_LUT4 C18141(
      .ADR0 (VCC),
      .ADR1 (syn24500),
      .ADR2 (VCC),
      .ADR3 (\bridge/conf_wb_img_ctrl1_out [1]),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/GROM )
    );
    X_INV \bridge/wishbone_slave_unit/wishbone_slave/mrl_en/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/wishbone_slave/mrl_en/YUSED (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/GROM ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/n_850 )
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/pref_en_reg (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/pref_en )
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/mrl_en/FFY/ASYNC_FF_GSR_OR_319 (
      .I0 (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/wishbone_slave/mrl_en_reg (
      .I (\bridge/wishbone_slave_unit/wishbone_slave/n_850 ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/wishbone_slave/C77/N9 ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en )
    );
    X_OR2
     \bridge/wishbone_slave_unit/wishbone_slave/mrl_en/FFX/ASYNC_FF_GSR_OR_320 (
      .I0 (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/wishbone_slave/mrl_en/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C17816.INIT = 16'hF0AA;
    X_LUT4 C17816(
      .ADR0 (\bridge/pci_target_unit/wishbone_master/N3116 ),
      .ADR1 (VCC),
      .ADR2 (\bridge/conf_cache_line_size_out [6]),
      .ADR3 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .O (\bridge/pci_target_unit/wishbone_master/C3414/N42 )
    );
    defparam C17815.INIT = 16'hACAC;
    X_LUT4 C17815(
      .ADR0 (\bridge/conf_cache_line_size_out [7]),
      .ADR1 (\bridge/pci_target_unit/wishbone_master/N3117 ),
      .ADR2 (\bridge/pci_target_unit/wishbone_master/C82/C0 ),
      .ADR3 (VCC),
      .O (\bridge/pci_target_unit/wishbone_master/C3414/N48 )
    );
    X_INV \bridge/pci_target_unit/wishbone_master/cache_line<7>/SRMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line[7]/SRNOT )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/cache_line_reg<6> (
      .I (\bridge/pci_target_unit/wishbone_master/C3414/N42 ),
      .CLK (CLK_BUFGPed),
      .CE (N12510),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/cache_line[7]/FFY/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line [6])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/cache_line<7>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/cache_line[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/cache_line[7]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/pci_target_unit/wishbone_master/cache_line_reg<7> (
      .I (\bridge/pci_target_unit/wishbone_master/C3414/N48 ),
      .CLK (CLK_BUFGPed),
      .CE (N12510),
      .SET (GND),
      .RST 
      (\bridge/pci_target_unit/wishbone_master/cache_line[7]/FFX/ASYNC_FF_GSR_OR ),
      .O (\bridge/pci_target_unit/wishbone_master/cache_line [7])
    );
    X_OR2
     \bridge/pci_target_unit/wishbone_master/cache_line<7>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/pci_target_unit/wishbone_master/cache_line[7]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/pci_target_unit/wishbone_master/cache_line[7]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam C18196.INIT = 16'h33CC;
    X_LUT4 C18196(
      .ADR0 (VCC),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [0]),
      .ADR2 (VCC),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [1]),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/GROM )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/SRNOT )
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<1>/YUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/GROM ),
      .O (\bridge/wishbone_slave_unit/fifos/outNextGreyCount [0])
    );
    X_FF \bridge/wishbone_slave_unit/fifos/outGreyCount_reg<0> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/GROM ),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/FFY/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/outGreyCount [0])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/FFY/ASYNC_FF_GSR_OR )

    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/outNextGreyCount [0]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/out_count_en ),
      .SET (GND),
      .RST 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/FFX/ASYNC_FF_GSR_OR )
,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount<1>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount[1]/FFX/ASYNC_FF_GSR_OR )

    );
    defparam C17749.INIT = 16'h00F0;
    X_LUT4 C17749(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty ),
      .ADR3 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/wclock_nempty_detect ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty111 )
    );
    defparam C19400.INIT = 16'h000A;
    X_LUT4 C19400(
      .ADR0 (syn19088),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/empty ),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty ),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/FROM )
    );
    X_INV
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/SRMUX (
      .I (N_RST),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/SRNOT )
    );
    X_BUF
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/XUSED (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/FROM )
      ,
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/rallow_out )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty_reg (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty111 ),
      .CLK (CLK_BUFGPed),
      .CE (VCC),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR )
,
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty )
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR_321 (
      .I0 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/wbw_fifo_ctrl/stretched_empty/FFY/ASYNC_FF_GSR_OR )

    );
    defparam C18197.INIT = 16'h0FF0;
    X_LUT4 C18197(
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [2]),
      .ADR3 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [1]),
      .O (\bridge/wishbone_slave_unit/fifos/outNextGreyCount [1])
    );
    X_INV \bridge/wishbone_slave_unit/fifos/outGreyCount<1>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/outGreyCount[1]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/outGreyCount_reg<1> (
      .I (\bridge/wishbone_slave_unit/fifos/outNextGreyCount [1]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/out_count_en ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/outGreyCount[1]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/outGreyCount [1])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/outGreyCount<1>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/outGreyCount[1]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/outGreyCount[1]/FFY/ASYNC_FF_GSR_OR )
    );
    defparam C18195.INIT = 16'h6666;
    X_LUT4 C18195(
      .ADR0 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [3]),
      .ADR1 (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [2]),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (\bridge/wishbone_slave_unit/fifos/outNextGreyCount [2])
    );
    X_INV \bridge/wishbone_slave_unit/fifos/outGreyCount<3>/SRMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/outGreyCount[3]/SRNOT )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/outGreyCount_reg<2> (
      .I (\bridge/wishbone_slave_unit/fifos/outNextGreyCount [2]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/out_count_en ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/outGreyCount[3]/FFY/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/outGreyCount [2])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/outGreyCount<3>/FFY/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/outGreyCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/outGreyCount[3]/FFY/ASYNC_FF_GSR_OR )
    );
    X_FF \bridge/wishbone_slave_unit/fifos/outGreyCount_reg<3> (
      .I (\bridge/wishbone_slave_unit/fifos/wbw_outTransactionCount [3]),
      .CLK (CLK_BUFGPed),
      .CE (\bridge/wishbone_slave_unit/fifos/out_count_en ),
      .SET 
      (\bridge/wishbone_slave_unit/fifos/outGreyCount[3]/FFX/ASYNC_FF_GSR_OR ),
      .RST (GND),
      .O (\bridge/wishbone_slave_unit/fifos/outGreyCount [3])
    );
    X_OR2
     \bridge/wishbone_slave_unit/fifos/outGreyCount<3>/FFX/ASYNC_FF_GSR_OR (
      .I0 (\bridge/wishbone_slave_unit/fifos/outGreyCount[3]/SRNOT ),
      .I1 (GSR),
      .O 
      (\bridge/wishbone_slave_unit/fifos/outGreyCount[3]/FFX/ASYNC_FF_GSR_OR )
    );
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_1 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S16_S16 \bridge/wishbone_slave_unit/fifos/dpram16_1 (
      .CLKA (CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\bridge/wishbone_slave_unit/fifos/dpram16_1/LOGIC_ONE ),
      .ENB (\bridge/wishbone_slave_unit/fifos/dpram16_1/LOGIC_ONE ),
      .RSTA (\bridge/wishbone_slave_unit/fifos/dpram16_1/RSTANOT ),
      .RSTB (\bridge/wishbone_slave_unit/fifos/dpram16_1/RSTBNOT ),
      .WEA (\bridge/wishbone_slave_unit/fifos/dpram16_1/WEANOT ),
      .WEB (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .GSR (GSR),
      .ADDRA ({N12607, N12607, \bridge/wishbone_slave_unit/fifos/C6/N35 , 
      \bridge/wishbone_slave_unit/fifos/C6/N30 , 
      \bridge/wishbone_slave_unit/fifos/C6/N24 , 
      \bridge/wishbone_slave_unit/fifos/C6/N18 , 
      \bridge/wishbone_slave_unit/fifos/C6/N12 , 
      \bridge/wishbone_slave_unit/fifos/C6/N6 }),
      .ADDRB ({\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out , 
      \bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out , 
      \bridge/wishbone_slave_unit/fifos/C3/N33 , 
      \bridge/wishbone_slave_unit/fifos/C3/N30 , 
      \bridge/wishbone_slave_unit/fifos/C3/N24 , 
      \bridge/wishbone_slave_unit/fifos/C3/N18 , 
      \bridge/wishbone_slave_unit/fifos/C3/N12 , 
      \bridge/wishbone_slave_unit/fifos/C3/N6 }),
      .DIA ({\bridge/wishbone_slave_unit/wbs_sm_data_out [15], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [14], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [13], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [12], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [11], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [10], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [9], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [8], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [7], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [6], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [5], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [4], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [3], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [2], GLOBAL_LOGIC0_7, 
      GLOBAL_LOGIC0_6}),
      .DIB ({\bridge/wishbone_slave_unit/pcim_sm_data_out [15], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [14], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [13], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [12], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [11], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [10], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [9], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [8], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [7], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [6], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [5], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [4], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [3], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [2], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [1], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [0]}),
      .DOA ({\bridge/wishbone_slave_unit/fifos_wbr_data_out [15], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [14], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [13], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [12], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [11], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [10], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [9], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [8], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [7], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [6], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [5], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [4], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [3], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [2], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [1], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [0]}),
      .DOB ({\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [15], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [14], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [13], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [12], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [11], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [10], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [9], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [8], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [7], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [6], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [5], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [4], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [3], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [2], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [1], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [0]})
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/dpram16_1/ANCHOR_PRIM (
      .I (\bridge/wishbone_slave_unit/fifos/dpram16_1/INT_SIG ),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_1/INT_SIG )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_1/WEAMUX (
      .I (N12607),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_1/WEANOT )
    );
    X_ONE \bridge/wishbone_slave_unit/fifos/dpram16_1/LOGIC_ONE_322 (
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_1/LOGIC_ONE )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_1/RSTAMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_1/RSTANOT )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_1/RSTBMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_1/RSTBNOT )
    );
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_2 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S16_S16 \bridge/wishbone_slave_unit/fifos/dpram16_2 (
      .CLKA (CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\bridge/wishbone_slave_unit/fifos/dpram16_2/LOGIC_ONE ),
      .ENB (\bridge/wishbone_slave_unit/fifos/dpram16_2/LOGIC_ONE ),
      .RSTA (\bridge/wishbone_slave_unit/fifos/dpram16_2/RSTANOT ),
      .RSTB (\bridge/wishbone_slave_unit/fifos/dpram16_2/RSTBNOT ),
      .WEA (\bridge/wishbone_slave_unit/fifos/dpram16_2/WEANOT ),
      .WEB (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .GSR (GSR),
      .ADDRA ({N12607, N12607, \bridge/wishbone_slave_unit/fifos/C6/N35 , 
      \bridge/wishbone_slave_unit/fifos/C6/N30 , 
      \bridge/wishbone_slave_unit/fifos/C6/N24 , 
      \bridge/wishbone_slave_unit/fifos/C6/N18 , 
      \bridge/wishbone_slave_unit/fifos/C6/N12 , 
      \bridge/wishbone_slave_unit/fifos/C6/N6 }),
      .ADDRB ({\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out , 
      \bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out , 
      \bridge/wishbone_slave_unit/fifos/C3/N33 , 
      \bridge/wishbone_slave_unit/fifos/C3/N30 , 
      \bridge/wishbone_slave_unit/fifos/C3/N24 , 
      \bridge/wishbone_slave_unit/fifos/C3/N18 , 
      \bridge/wishbone_slave_unit/fifos/C3/N12 , 
      \bridge/wishbone_slave_unit/fifos/C3/N6 }),
      .DIA ({\bridge/wishbone_slave_unit/wbs_sm_data_out [31], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [30], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [29], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [28], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [27], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [26], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [25], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [24], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [23], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [22], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [21], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [20], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [19], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [18], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [17], 
      \bridge/wishbone_slave_unit/wbs_sm_data_out [16]}),
      .DIB ({\bridge/wishbone_slave_unit/pcim_sm_data_out [31], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [30], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [29], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [28], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [27], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [26], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [25], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [24], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [23], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [22], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [21], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [20], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [19], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [18], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [17], 
      \bridge/wishbone_slave_unit/pcim_sm_data_out [16]}),
      .DOA ({\bridge/wishbone_slave_unit/fifos_wbr_data_out [31], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [30], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [29], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [28], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [27], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [26], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [25], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [24], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [23], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [22], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [21], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [20], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [19], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [18], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [17], 
      \bridge/wishbone_slave_unit/fifos_wbr_data_out [16]}),
      .DOB ({\bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [31], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [30], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [29], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [28], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [27], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [26], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [25], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [24], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [23], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [22], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [21], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [20], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [19], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [18], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [17], 
      \bridge/wishbone_slave_unit/fifos_wbw_addr_data_out [16]})
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/dpram16_2/ANCHOR_PRIM (
      .I (\bridge/wishbone_slave_unit/fifos/dpram16_2/INT_SIG ),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_2/INT_SIG )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_2/WEAMUX (
      .I (N12607),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_2/WEANOT )
    );
    X_ONE \bridge/wishbone_slave_unit/fifos/dpram16_2/LOGIC_ONE_323 (
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_2/LOGIC_ONE )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_2/RSTAMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_2/RSTANOT )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_2/RSTBMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_2/RSTBNOT )
    );
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/wishbone_slave_unit/fifos/dpram16_3 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S16_S16 \bridge/wishbone_slave_unit/fifos/dpram16_3 (
      .CLKA (CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\bridge/wishbone_slave_unit/fifos/dpram16_3/LOGIC_ONE ),
      .ENB (\bridge/wishbone_slave_unit/fifos/dpram16_3/LOGIC_ONE ),
      .RSTA (\bridge/wishbone_slave_unit/fifos/dpram16_3/RSTANOT ),
      .RSTB (\bridge/wishbone_slave_unit/fifos/dpram16_3/RSTBNOT ),
      .WEA (\bridge/wishbone_slave_unit/fifos/dpram16_3/WEANOT ),
      .WEB (\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out ),
      .GSR (GSR),
      .ADDRA ({N12607, N12607, \bridge/wishbone_slave_unit/fifos/C6/N35 , 
      \bridge/wishbone_slave_unit/fifos/C6/N30 , 
      \bridge/wishbone_slave_unit/fifos/C6/N24 , 
      \bridge/wishbone_slave_unit/fifos/C6/N18 , 
      \bridge/wishbone_slave_unit/fifos/C6/N12 , 
      \bridge/wishbone_slave_unit/fifos/C6/N6 }),
      .ADDRB ({\bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out , 
      \bridge/wishbone_slave_unit/pcim_if_wbr_wenable_out , 
      \bridge/wishbone_slave_unit/fifos/C3/N33 , 
      \bridge/wishbone_slave_unit/fifos/C3/N30 , 
      \bridge/wishbone_slave_unit/fifos/C3/N24 , 
      \bridge/wishbone_slave_unit/fifos/C3/N18 , 
      \bridge/wishbone_slave_unit/fifos/C3/N12 , 
      \bridge/wishbone_slave_unit/fifos/C3/N6 }),
      .DIA ({N12360, GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_9, 
      \bridge/wishbone_slave_unit/wbs_sm_wbw_control_out [0], GLOBAL_LOGIC0_11, 
      GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_11, GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_3, 
      GLOBAL_LOGIC0_8, GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_9, 
      \bridge/wishbone_slave_unit/wbs_sm_cbe_out [3], 
      \bridge/wishbone_slave_unit/wbs_sm_cbe_out [2], GLOBAL_LOGIC1, GLOBAL_LOGIC1}),
      .DIB ({GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_9, 
      \bridge/wishbone_slave_unit/pcim_if_wbr_control_out [1], 
      \bridge/wishbone_slave_unit/pcim_if_wbr_control_out [0], GLOBAL_LOGIC0_11, 
      GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_11, GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_9, 
      GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_9, 
      \bridge/wishbone_slave_unit/pcim_if_wbr_be_out [3], 
      \bridge/wishbone_slave_unit/pcim_if_wbr_be_out [2], 
      \bridge/wishbone_slave_unit/pcim_if_wbr_be_out [1], 
      \bridge/wishbone_slave_unit/pcim_if_wbr_be_out [0]}),
      .DOA ({\bridge/wishbone_slave_unit/fifos/dpram16_3/DOA15 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA14 , 
      \bridge/wishbone_slave_unit/fifos_wbr_control_out [1], 
      \bridge/wishbone_slave_unit/fifos_wbr_control_out [0], 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA11 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA10 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA9 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA8 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA7 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA6 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA5 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA4 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA3 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA2 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA1 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOA0 }),
      .DOB ({\bridge/wishbone_slave_unit/fifos/dpram16_3/DOB15 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB14 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB13 , 
      \bridge/wishbone_slave_unit/fifos_wbw_control_out [0], 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB11 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB10 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB9 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB8 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB7 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB6 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB5 , 
      \bridge/wishbone_slave_unit/fifos/dpram16_3/DOB4 , 
      \bridge/wishbone_slave_unit/fifos_wbw_cbe_out [3], 
      \bridge/wishbone_slave_unit/fifos_wbw_cbe_out [2], 
      \bridge/wishbone_slave_unit/fifos_wbw_cbe_out [1], 
      \bridge/wishbone_slave_unit/fifos_wbw_cbe_out [0]})
    );
    X_BUF \bridge/wishbone_slave_unit/fifos/dpram16_3/ANCHOR_PRIM (
      .I (\bridge/wishbone_slave_unit/fifos/dpram16_3/INT_SIG ),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_3/INT_SIG )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_3/WEAMUX (
      .I (N12607),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_3/WEANOT )
    );
    X_ONE \bridge/wishbone_slave_unit/fifos/dpram16_3/LOGIC_ONE_324 (
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_3/LOGIC_ONE )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_3/RSTAMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_3/RSTANOT )
    );
    X_INV \bridge/wishbone_slave_unit/fifos/dpram16_3/RSTBMUX (
      .I (N_RST),
      .O (\bridge/wishbone_slave_unit/fifos/dpram16_3/RSTBNOT )
    );
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_0 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S8_S16 \CRT/ssvga_fifo/ramb4_s8_0 (
      .CLKA (CRT_CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ONE ),
      .ENB (\CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ONE ),
      .RSTA (\CRT/ssvga_fifo/ramb4_s8_0/RSTANOT ),
      .RSTB (\CRT/ssvga_fifo/ramb4_s8_0/RSTBNOT ),
      .WEA (\CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ZERO ),
      .WEB (\CRT/fifo_wr_en ),
      .GSR (GSR),
      .ADDRA ({\CRT/ssvga_fifo/C6/N54 , \CRT/ssvga_fifo/C6/N48 , 
      \CRT/ssvga_fifo/C6/N42 , \CRT/ssvga_fifo/C6/N36 , \CRT/ssvga_fifo/C6/N30 , 
      \CRT/ssvga_fifo/C6/N24 , \CRT/ssvga_fifo/C6/N18 , \CRT/ssvga_fifo/C6/N12 , 
      \CRT/ssvga_fifo/C6/N6 }),
      .ADDRB ({\CRT/ssvga_fifo/wr_ptr [7], \CRT/ssvga_fifo/wr_ptr [6], 
      \CRT/ssvga_fifo/wr_ptr [5], \CRT/ssvga_fifo/wr_ptr [4], 
      \CRT/ssvga_fifo/wr_ptr [3], \CRT/ssvga_fifo/wr_ptr [2], 
      \CRT/ssvga_fifo/wr_ptr [1], \CRT/ssvga_fifo/wr_ptr [0]}),
      .DIA ({GLOBAL_LOGIC0_2, GLOBAL_LOGIC0_2, GLOBAL_LOGIC0_1, GLOBAL_LOGIC0_1
      , GLOBAL_LOGIC0_1, GLOBAL_LOGIC0_2, GLOBAL_LOGIC0_1, GLOBAL_LOGIC0_2}),
      .DIB ({SDAT_O[15], SDAT_O[14], SDAT_O[13], SDAT_O[12], SDAT_O[11], 
      SDAT_O[10], SDAT_O[9], SDAT_O[8], SDAT_O[7], SDAT_O[6], SDAT_O[5], SDAT_O[4], 
      SDAT_O[3], SDAT_O[2], SDAT_O[1], SDAT_O[0]}),
      .DOA ({\CRT/ssvga_fifo/dat_o_low [7], \CRT/ssvga_fifo/dat_o_low [6], 
      \CRT/ssvga_fifo/dat_o_low [5], \CRT/ssvga_fifo/dat_o_low [4], 
      \CRT/ssvga_fifo/dat_o_low [3], \CRT/ssvga_fifo/dat_o_low [2], 
      \CRT/ssvga_fifo/dat_o_low [1], \CRT/ssvga_fifo/dat_o_low [0]}),
      .DOB ({\CRT/ssvga_fifo/ramb4_s8_0/DOB15 , 
      \CRT/ssvga_fifo/ramb4_s8_0/DOB14 , \CRT/ssvga_fifo/ramb4_s8_0/DOB13 , 
      \CRT/ssvga_fifo/ramb4_s8_0/DOB12 , \CRT/ssvga_fifo/ramb4_s8_0/DOB11 , 
      \CRT/ssvga_fifo/ramb4_s8_0/DOB10 , \CRT/ssvga_fifo/ramb4_s8_0/DOB9 , 
      \CRT/ssvga_fifo/ramb4_s8_0/DOB8 , \CRT/ssvga_fifo/ramb4_s8_0/DOB7 , 
      \CRT/ssvga_fifo/ramb4_s8_0/DOB6 , \CRT/ssvga_fifo/ramb4_s8_0/DOB5 , 
      \CRT/ssvga_fifo/ramb4_s8_0/DOB4 , \CRT/ssvga_fifo/ramb4_s8_0/DOB3 , 
      \CRT/ssvga_fifo/ramb4_s8_0/DOB2 , \CRT/ssvga_fifo/ramb4_s8_0/DOB1 , 
      \CRT/ssvga_fifo/ramb4_s8_0/DOB0 })
    );
    X_BUF \CRT/ssvga_fifo/ramb4_s8_0/ANCHOR_PRIM (
      .I (\CRT/ssvga_fifo/ramb4_s8_0/INT_SIG ),
      .O (\CRT/ssvga_fifo/ramb4_s8_0/INT_SIG )
    );
    X_ZERO \CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ZERO_325 (
      .O (\CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ZERO )
    );
    X_ONE \CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ONE_326 (
      .O (\CRT/ssvga_fifo/ramb4_s8_0/LOGIC_ONE )
    );
    X_INV \CRT/ssvga_fifo/ramb4_s8_0/RSTAMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/ramb4_s8_0/RSTANOT )
    );
    X_INV \CRT/ssvga_fifo/ramb4_s8_0/RSTBMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/ramb4_s8_0/RSTBNOT )
    );
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_fifo/ramb4_s8_1 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S8_S16 \CRT/ssvga_fifo/ramb4_s8_1 (
      .CLKA (CRT_CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ONE ),
      .ENB (\CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ONE ),
      .RSTA (\CRT/ssvga_fifo/ramb4_s8_1/RSTANOT ),
      .RSTB (\CRT/ssvga_fifo/ramb4_s8_1/RSTBNOT ),
      .WEA (\CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ZERO ),
      .WEB (\CRT/fifo_wr_en ),
      .GSR (GSR),
      .ADDRA ({\CRT/ssvga_fifo/C6/N54 , \CRT/ssvga_fifo/C6/N48 , 
      \CRT/ssvga_fifo/C6/N42 , \CRT/ssvga_fifo/C6/N36 , \CRT/ssvga_fifo/C6/N30 , 
      \CRT/ssvga_fifo/C6/N24 , \CRT/ssvga_fifo/C6/N18 , \CRT/ssvga_fifo/C6/N12 , 
      \CRT/ssvga_fifo/C6/N6 }),
      .ADDRB ({\CRT/ssvga_fifo/wr_ptr [7], \CRT/ssvga_fifo/wr_ptr [6], 
      \CRT/ssvga_fifo/wr_ptr [5], \CRT/ssvga_fifo/wr_ptr [4], 
      \CRT/ssvga_fifo/wr_ptr [3], \CRT/ssvga_fifo/wr_ptr [2], 
      \CRT/ssvga_fifo/wr_ptr [1], \CRT/ssvga_fifo/wr_ptr [0]}),
      .DIA ({GLOBAL_LOGIC0_8, GLOBAL_LOGIC0_8, GLOBAL_LOGIC0_9, GLOBAL_LOGIC0_8
      , GLOBAL_LOGIC0_10, GLOBAL_LOGIC0_8, GLOBAL_LOGIC0_10, GLOBAL_LOGIC0_8}),
      .DIB ({SDAT_O[31], SDAT_O[30], SDAT_O[29], SDAT_O[28], SDAT_O[27], 
      SDAT_O[26], SDAT_O[25], SDAT_O[24], SDAT_O[23], SDAT_O[22], SDAT_O[21], 
      SDAT_O[20], SDAT_O[19], SDAT_O[18], SDAT_O[17], SDAT_O[16]}),
      .DOA ({\CRT/ssvga_fifo/dat_o_high [7], \CRT/ssvga_fifo/dat_o_high [6], 
      \CRT/ssvga_fifo/dat_o_high [5], \CRT/ssvga_fifo/dat_o_high [4], 
      \CRT/ssvga_fifo/dat_o_high [3], \CRT/ssvga_fifo/dat_o_high [2], 
      \CRT/ssvga_fifo/dat_o_high [1], \CRT/ssvga_fifo/dat_o_high [0]}),
      .DOB ({\CRT/ssvga_fifo/ramb4_s8_1/DOB15 , 
      \CRT/ssvga_fifo/ramb4_s8_1/DOB14 , \CRT/ssvga_fifo/ramb4_s8_1/DOB13 , 
      \CRT/ssvga_fifo/ramb4_s8_1/DOB12 , \CRT/ssvga_fifo/ramb4_s8_1/DOB11 , 
      \CRT/ssvga_fifo/ramb4_s8_1/DOB10 , \CRT/ssvga_fifo/ramb4_s8_1/DOB9 , 
      \CRT/ssvga_fifo/ramb4_s8_1/DOB8 , \CRT/ssvga_fifo/ramb4_s8_1/DOB7 , 
      \CRT/ssvga_fifo/ramb4_s8_1/DOB6 , \CRT/ssvga_fifo/ramb4_s8_1/DOB5 , 
      \CRT/ssvga_fifo/ramb4_s8_1/DOB4 , \CRT/ssvga_fifo/ramb4_s8_1/DOB3 , 
      \CRT/ssvga_fifo/ramb4_s8_1/DOB2 , \CRT/ssvga_fifo/ramb4_s8_1/DOB1 , 
      \CRT/ssvga_fifo/ramb4_s8_1/DOB0 })
    );
    X_BUF \CRT/ssvga_fifo/ramb4_s8_1/ANCHOR_PRIM (
      .I (\CRT/ssvga_fifo/ramb4_s8_1/INT_SIG ),
      .O (\CRT/ssvga_fifo/ramb4_s8_1/INT_SIG )
    );
    X_ZERO \CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ZERO_327 (
      .O (\CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ZERO )
    );
    X_ONE \CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ONE_328 (
      .O (\CRT/ssvga_fifo/ramb4_s8_1/LOGIC_ONE )
    );
    X_INV \CRT/ssvga_fifo/ramb4_s8_1/RSTAMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/ramb4_s8_1/RSTANOT )
    );
    X_INV \CRT/ssvga_fifo/ramb4_s8_1/RSTBMUX (
      .I (N_RST),
      .O (\CRT/ssvga_fifo/ramb4_s8_1/RSTBNOT )
    );
    defparam \CRT/ssvga_pallete .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \CRT/ssvga_pallete .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S16_S16 \CRT/ssvga_pallete (
      .CLKA (CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\CRT/ssvga_pallete/LOGIC_ONE ),
      .ENB (\CRT/ssvga_pallete/LOGIC_ONE ),
      .RSTA (\CRT/ssvga_pallete/RSTANOT ),
      .RSTB (\CRT/ssvga_pallete/RSTBNOT ),
      .WEA (\CRT/pal_wr_en ),
      .WEB (\CRT/ssvga_pallete/LOGIC_ZERO ),
      .GSR (GSR),
      .ADDRA ({ADR_O[9], ADR_O[8], ADR_O[7], ADR_O[6], ADR_O[5], ADR_O[4], 
      ADR_O[3], ADR_O[2]}),
      .ADDRB ({\CRT/fifo_out [7], \CRT/fifo_out [6], \CRT/fifo_out [5], 
      \CRT/fifo_out [4], \CRT/fifo_out [3], \CRT/fifo_out [2], \CRT/fifo_out [1], 
      \CRT/fifo_out [0]}),
      .DIA ({\bridge/pci_target_unit/fifos_pciw_addr_data_out [15], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [14], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [13], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [12], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [11], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [10], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [9], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [8], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [7], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [6], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [5], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [4], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [3], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [2], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [1], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [0]}),
      .DIB ({GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_5, GLOBAL_LOGIC0_5
      , GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_5, GLOBAL_LOGIC0_5, GLOBAL_LOGIC0_5, 
      GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_5, GLOBAL_LOGIC0_4, 
      GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4, GLOBAL_LOGIC0_4}),
      .DOA ({\CRT/wbs_pal_data [15], \CRT/wbs_pal_data [14], 
      \CRT/wbs_pal_data [13], \CRT/wbs_pal_data [12], \CRT/wbs_pal_data [11], 
      \CRT/wbs_pal_data [10], \CRT/wbs_pal_data [9], \CRT/wbs_pal_data [8], 
      \CRT/wbs_pal_data [7], \CRT/wbs_pal_data [6], \CRT/wbs_pal_data [5], 
      \CRT/wbs_pal_data [4], \CRT/wbs_pal_data [3], \CRT/wbs_pal_data [2], 
      \CRT/wbs_pal_data [1], \CRT/wbs_pal_data [0]}),
      .DOB ({\CRT/pal_pix_dat [15], \CRT/pal_pix_dat [14], \CRT/pal_pix_dat [13]
      , \CRT/pal_pix_dat [12], \CRT/pal_pix_dat [11], \CRT/pal_pix_dat [10], 
      \CRT/pal_pix_dat [9], \CRT/pal_pix_dat [8], \CRT/pal_pix_dat [7], 
      \CRT/pal_pix_dat [6], \CRT/pal_pix_dat [5], \CRT/pal_pix_dat [4], 
      \CRT/ssvga_pallete/DOB3 , \CRT/ssvga_pallete/DOB2 , \CRT/ssvga_pallete/DOB1 , 
      \CRT/ssvga_pallete/DOB0 })
    );
    X_BUF \CRT/ssvga_pallete/ANCHOR_PRIM (
      .I (\CRT/ssvga_pallete/INT_SIG ),
      .O (\CRT/ssvga_pallete/INT_SIG )
    );
    X_ZERO \CRT/ssvga_pallete/LOGIC_ZERO_329 (
      .O (\CRT/ssvga_pallete/LOGIC_ZERO )
    );
    X_ONE \CRT/ssvga_pallete/LOGIC_ONE_330 (
      .O (\CRT/ssvga_pallete/LOGIC_ONE )
    );
    X_INV \CRT/ssvga_pallete/RSTAMUX (
      .I (N_RST),
      .O (\CRT/ssvga_pallete/RSTANOT )
    );
    X_INV \CRT/ssvga_pallete/RSTBMUX (
      .I (N_RST),
      .O (\CRT/ssvga_pallete/RSTBNOT )
    );
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_1 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S16_S16 \bridge/pci_target_unit/fifos/dpram16_1 (
      .CLKA (CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\bridge/pci_target_unit/fifos/portA_enable ),
      .ENB (\bridge/pci_target_unit/fifos/portB_enable ),
      .RSTA (\bridge/pci_target_unit/fifos/dpram16_1/RSTANOT ),
      .RSTB (\bridge/pci_target_unit/fifos/dpram16_1/RSTBNOT ),
      .WEA (\bridge/pci_target_unit/fifos/dpram16_1/WEANOT ),
      .WEB (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .GSR (GSR),
      .ADDRA ({N12616, N12616, N12616, \bridge/pci_target_unit/fifos/C9/N30 , 
      \bridge/pci_target_unit/fifos/C9/N24 , \bridge/pci_target_unit/fifos/C9/N18 , 
      \bridge/pci_target_unit/fifos/C9/N12 , \bridge/pci_target_unit/fifos/C9/N6 }),
      .ADDRB ({\bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/C10/N30 , \bridge/pci_target_unit/fifos/C10/N24 , 
      \bridge/pci_target_unit/fifos/C10/N18 , \bridge/pci_target_unit/fifos/C10/N12 , 
      \bridge/pci_target_unit/fifos/C10/N6 }),
      .DIA ({\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [15], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [14], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [13], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [12], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [11], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [10], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [9], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [8], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [7], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [6], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [5], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [4], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [3], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [2], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [1], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [0]}),
      .DIB ({\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [15], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [14], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [13], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [12], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [11], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [10], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [9], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [8], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [7], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [6], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [5], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [4], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [3], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [2], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [1], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [0]}),
      .DOA ({\bridge/pci_target_unit/fifos_pcir_data_out [15], 
      \bridge/pci_target_unit/fifos_pcir_data_out [14], 
      \bridge/pci_target_unit/fifos_pcir_data_out [13], 
      \bridge/pci_target_unit/fifos_pcir_data_out [12], 
      \bridge/pci_target_unit/fifos_pcir_data_out [11], 
      \bridge/pci_target_unit/fifos_pcir_data_out [10], 
      \bridge/pci_target_unit/fifos_pcir_data_out [9], 
      \bridge/pci_target_unit/fifos_pcir_data_out [8], 
      \bridge/pci_target_unit/fifos_pcir_data_out [7], 
      \bridge/pci_target_unit/fifos_pcir_data_out [6], 
      \bridge/pci_target_unit/fifos_pcir_data_out [5], 
      \bridge/pci_target_unit/fifos_pcir_data_out [4], 
      \bridge/pci_target_unit/fifos_pcir_data_out [3], 
      \bridge/pci_target_unit/fifos_pcir_data_out [2], 
      \bridge/pci_target_unit/fifos_pcir_data_out [1], 
      \bridge/pci_target_unit/fifos_pcir_data_out [0]}),
      .DOB ({\bridge/pci_target_unit/fifos_pciw_addr_data_out [15], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [14], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [13], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [12], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [11], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [10], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [9], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [8], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [7], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [6], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [5], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [4], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [3], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [2], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [1], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [0]})
    );
    X_BUF \bridge/pci_target_unit/fifos/dpram16_1/ANCHOR_PRIM (
      .I (\bridge/pci_target_unit/fifos/dpram16_1/INT_SIG ),
      .O (\bridge/pci_target_unit/fifos/dpram16_1/INT_SIG )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_1/WEAMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/dpram16_1/WEANOT )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_1/RSTAMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/dpram16_1/RSTANOT )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_1/RSTBMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/dpram16_1/RSTBNOT )
    );
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_2 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S16_S16 \bridge/pci_target_unit/fifos/dpram16_2 (
      .CLKA (CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\bridge/pci_target_unit/fifos/portA_enable ),
      .ENB (\bridge/pci_target_unit/fifos/portB_enable ),
      .RSTA (\bridge/pci_target_unit/fifos/dpram16_2/RSTANOT ),
      .RSTB (\bridge/pci_target_unit/fifos/dpram16_2/RSTBNOT ),
      .WEA (\bridge/pci_target_unit/fifos/dpram16_2/WEANOT ),
      .WEB (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .GSR (GSR),
      .ADDRA ({N12616, N12616, N12616, \bridge/pci_target_unit/fifos/C9/N30 , 
      \bridge/pci_target_unit/fifos/C9/N24 , \bridge/pci_target_unit/fifos/C9/N18 , 
      \bridge/pci_target_unit/fifos/C9/N12 , \bridge/pci_target_unit/fifos/C9/N6 }),
      .ADDRB ({\bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/C10/N30 , \bridge/pci_target_unit/fifos/C10/N24 , 
      \bridge/pci_target_unit/fifos/C10/N18 , \bridge/pci_target_unit/fifos/C10/N12 , 
      \bridge/pci_target_unit/fifos/C10/N6 }),
      .DIA ({\bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [31], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [30], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [29], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [28], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [27], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [26], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [25], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [24], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [23], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [22], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [21], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [20], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [19], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [18], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [17], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_addr_data_out [16]}),
      .DIB ({\bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [31], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [30], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [29], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [28], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [27], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [26], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [25], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [24], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [23], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [22], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [21], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [20], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [19], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [18], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [17], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_data_out [16]}),
      .DOA ({\bridge/pci_target_unit/fifos_pcir_data_out [31], 
      \bridge/pci_target_unit/fifos_pcir_data_out [30], 
      \bridge/pci_target_unit/fifos_pcir_data_out [29], 
      \bridge/pci_target_unit/fifos_pcir_data_out [28], 
      \bridge/pci_target_unit/fifos_pcir_data_out [27], 
      \bridge/pci_target_unit/fifos_pcir_data_out [26], 
      \bridge/pci_target_unit/fifos_pcir_data_out [25], 
      \bridge/pci_target_unit/fifos_pcir_data_out [24], 
      \bridge/pci_target_unit/fifos_pcir_data_out [23], 
      \bridge/pci_target_unit/fifos_pcir_data_out [22], 
      \bridge/pci_target_unit/fifos_pcir_data_out [21], 
      \bridge/pci_target_unit/fifos_pcir_data_out [20], 
      \bridge/pci_target_unit/fifos_pcir_data_out [19], 
      \bridge/pci_target_unit/fifos_pcir_data_out [18], 
      \bridge/pci_target_unit/fifos_pcir_data_out [17], 
      \bridge/pci_target_unit/fifos_pcir_data_out [16]}),
      .DOB ({\bridge/pci_target_unit/fifos_pciw_addr_data_out [31], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [30], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [29], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [28], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [27], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [26], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [25], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [24], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [23], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [22], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [21], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [20], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [19], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [18], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [17], 
      \bridge/pci_target_unit/fifos_pciw_addr_data_out [16]})
    );
    X_BUF \bridge/pci_target_unit/fifos/dpram16_2/ANCHOR_PRIM (
      .I (\bridge/pci_target_unit/fifos/dpram16_2/INT_SIG ),
      .O (\bridge/pci_target_unit/fifos/dpram16_2/INT_SIG )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_2/WEAMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/dpram16_2/WEANOT )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_2/RSTAMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/dpram16_2/RSTANOT )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_2/RSTBMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/dpram16_2/RSTBNOT )
    );
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \bridge/pci_target_unit/fifos/dpram16_3 .INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    X_RAMB4_S16_S16 \bridge/pci_target_unit/fifos/dpram16_3 (
      .CLKA (CLK_BUFGPed),
      .CLKB (CLK_BUFGPed),
      .ENA (\bridge/pci_target_unit/fifos/portA_enable ),
      .ENB (\bridge/pci_target_unit/fifos/portB_enable ),
      .RSTA (\bridge/pci_target_unit/fifos/dpram16_3/RSTANOT ),
      .RSTB (\bridge/pci_target_unit/fifos/dpram16_3/RSTBNOT ),
      .WEA (\bridge/pci_target_unit/fifos/dpram16_3/WEANOT ),
      .WEB (\bridge/pci_target_unit/fifos/pcir_wallow ),
      .GSR (GSR),
      .ADDRA ({N12616, N12616, N12616, \bridge/pci_target_unit/fifos/C9/N30 , 
      \bridge/pci_target_unit/fifos/C9/N24 , \bridge/pci_target_unit/fifos/C9/N18 , 
      \bridge/pci_target_unit/fifos/C9/N12 , \bridge/pci_target_unit/fifos/C9/N6 }),
      .ADDRB ({\bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/pcir_wallow , 
      \bridge/pci_target_unit/fifos/C10/N30 , \bridge/pci_target_unit/fifos/C10/N24 , 
      \bridge/pci_target_unit/fifos/C10/N18 , \bridge/pci_target_unit/fifos/C10/N12 , 
      \bridge/pci_target_unit/fifos/C10/N6 }),
      .DIA ({GLOBAL_LOGIC0_0, 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_control_out[2] , GLOBAL_LOGIC0, 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_control_out[0] , GLOBAL_LOGIC0, 
      GLOBAL_LOGIC0_0, GLOBAL_LOGIC0, GLOBAL_LOGIC0, GLOBAL_LOGIC0, GLOBAL_LOGIC0, 
      GLOBAL_LOGIC0, GLOBAL_LOGIC0, 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out [3], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out [2], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out [1], 
      \bridge/pci_target_unit/pcit_if_pciw_fifo_cbe_out [0]}),
      .DIB ({GLOBAL_LOGIC0_0, GLOBAL_LOGIC0_0, 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out [1], 
      \bridge/pci_target_unit/wbm_sm_pcir_fifo_control_out [0], GLOBAL_LOGIC0_0, 
      GLOBAL_LOGIC0, GLOBAL_LOGIC0_0, GLOBAL_LOGIC0, GLOBAL_LOGIC0_0, GLOBAL_LOGIC0_0
      , GLOBAL_LOGIC0, GLOBAL_LOGIC0, \bridge/pci_target_unit/del_sync_be_out [3], 
      \bridge/pci_target_unit/del_sync_be_out [2], 
      \bridge/pci_target_unit/del_sync_be_out [1], 
      \bridge/pci_target_unit/del_sync_be_out [0]}),
      .DOA ({\bridge/pci_target_unit/fifos/dpram16_3/DOA15 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA14 , 
      \bridge/pci_target_unit/fifos_pcir_control_out [1], 
      \bridge/pci_target_unit/fifos_pcir_control_out [0], 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA11 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA10 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA9 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA8 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA7 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA6 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA5 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA4 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA3 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA2 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA1 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOA0 }),
      .DOB ({\bridge/pci_target_unit/fifos/dpram16_3/DOB15 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB14 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB13 , 
      \bridge/pci_target_unit/fifos_pciw_control_out [0], 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB11 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB10 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB9 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB8 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB7 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB6 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB5 , 
      \bridge/pci_target_unit/fifos/dpram16_3/DOB4 , 
      \bridge/pci_target_unit/fifos_pciw_cbe_out [3], 
      \bridge/pci_target_unit/fifos_pciw_cbe_out [2], 
      \bridge/pci_target_unit/fifos_pciw_cbe_out [1], 
      \bridge/pci_target_unit/fifos_pciw_cbe_out [0]})
    );
    X_BUF \bridge/pci_target_unit/fifos/dpram16_3/ANCHOR_PRIM (
      .I (\bridge/pci_target_unit/fifos/dpram16_3/INT_SIG ),
      .O (\bridge/pci_target_unit/fifos/dpram16_3/INT_SIG )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_3/WEAMUX (
      .I (N12616),
      .O (\bridge/pci_target_unit/fifos/dpram16_3/WEANOT )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_3/RSTAMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/dpram16_3/RSTANOT )
    );
    X_INV \bridge/pci_target_unit/fifos/dpram16_3/RSTBMUX (
      .I (N_RST),
      .O (\bridge/pci_target_unit/fifos/dpram16_3/RSTBNOT )
    );
    X_CKBUF \CLK/BUF (
      .I (CLK),
      .O (\C20042/IBUFG )
    );
    X_IPAD \CLK/PAD (
      .PAD (CLK)
    );
    X_CKBUF \CRT_CLK/BUF (
      .I (CRT_CLK),
      .O (\C20043/IBUFG )
    );
    X_IPAD \CRT_CLK/PAD (
      .PAD (CRT_CLK)
    );
    X_CKBUF \C20042/BUFG/BUF (
      .I (\C20042/IBUFG ),
      .O (CLK_BUFGPed)
    );
    X_CKBUF \C20043/BUFG/BUF (
      .I (\C20043/IBUFG ),
      .O (CRT_CLK_BUFGPed)
    );
    defparam \PWR_GND_0/G .INIT = 16'h0000;
    X_LUT4 \PWR_GND_0/G (
      .ADR0 (VCC),
      .ADR1 (VCC),
      .ADR2 (VCC),
      .ADR3 (VCC),
      .O (GLOBAL_LOGIC0_10)
    );
    X_INV \AD<27>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[27]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<26>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[26]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<25>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[25]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<24>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[24]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<23>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[23]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \CBE<3>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\CBE[3]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<17>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[17]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<16>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[16]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \CBE<2>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\CBE[2]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \STOP/OUTBUF_GTS_AND_1_INV_331 (
      .I (GTS),
      .O (\STOP/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<22>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[22]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \FRAME/OUTBUF_GTS_AND_1_INV_332 (
      .I (GTS),
      .O (\FRAME/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \PERR/OUTBUF_GTS_AND_1_INV_333 (
      .I (GTS),
      .O (\PERR/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<21>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[21]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \IRDY/OUTBUF_GTS_AND_1_INV_334 (
      .I (GTS),
      .O (\IRDY/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<20>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[20]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \SERR/OUTBUF_GTS_AND_1_INV_335 (
      .I (GTS),
      .O (\SERR/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<19>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[19]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<13>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[13]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \PAR/OUTBUF_GTS_AND_1_INV_336 (
      .I (GTS),
      .O (\PAR/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<18>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[18]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<12>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[12]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \CBE<1>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\CBE[1]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \TRDY/OUTBUF_GTS_AND_1_INV_337 (
      .I (GTS),
      .O (\TRDY/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<11>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[11]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<15>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[15]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<14>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[14]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \DEVSEL/OUTBUF_GTS_AND_1_INV_338 (
      .I (GTS),
      .O (\DEVSEL/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<10>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[10]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<3>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[3]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<9>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[9]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<2>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[2]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<8>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[8]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<1>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[1]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \CBE<0>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\CBE[0]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<6>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[6]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<7>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[7]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<5>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[5]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV C_HSYNC_2_INV_339(
      .I (GTS),
      .O (C_HSYNC_2_INV)
    );
    X_INV \AD<4>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[4]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \REQ/OUTBUF_GTS_AND_1_INV_340 (
      .I (GTS),
      .O (\REQ/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<0>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[0]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV C_VSYNC_2_INV_341(
      .I (GTS),
      .O (C_VSYNC_2_INV)
    );
    X_INV C_LED_2_INV_342(
      .I (GTS),
      .O (C_LED_2_INV)
    );
    X_INV \AD<31>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[31]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<30>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[30]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<29>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[29]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \AD<28>/OUTBUF_GTS_AND_1_INV (
      .I (GTS),
      .O (\AD[28]/OUTBUF_GTS_AND_1_INV )
    );
    X_INV \C_RGB<14>_2_INV (
      .I (GTS),
      .O (\C_RGB[14]_2_INV )
    );
    X_INV \C_RGB<7>_2_INV (
      .I (GTS),
      .O (\C_RGB[7]_2_INV )
    );
    X_INV \C_RGB<15>_2_INV (
      .I (GTS),
      .O (\C_RGB[15]_2_INV )
    );
    X_INV \C_RGB<8>_2_INV (
      .I (GTS),
      .O (\C_RGB[8]_2_INV )
    );
    X_INV \C_RGB<9>_2_INV (
      .I (GTS),
      .O (\C_RGB[9]_2_INV )
    );
    X_INV \C_RGB<4>_2_INV (
      .I (GTS),
      .O (\C_RGB[4]_2_INV )
    );
    X_INV \C_RGB<5>_2_INV (
      .I (GTS),
      .O (\C_RGB[5]_2_INV )
    );
    X_INV \C_RGB<10>_2_INV (
      .I (GTS),
      .O (\C_RGB[10]_2_INV )
    );
    X_INV \C_RGB<6>_2_INV (
      .I (GTS),
      .O (\C_RGB[6]_2_INV )
    );
    X_INV \C_RGB<11>_2_INV (
      .I (GTS),
      .O (\C_RGB[11]_2_INV )
    );
    X_INV \C_RGB<12>_2_INV (
      .I (GTS),
      .O (\C_RGB[12]_2_INV )
    );
    X_INV \C_RGB<13>_2_INV (
      .I (GTS),
      .O (\C_RGB[13]_2_INV )
    );
    X_ONE VCC_343(
      .O (VCC)
    );
    X_ZERO GND_344(
      .O (GND)
    );
    X_PD NGD2VER_PD_9881 (.O (GSR) );
    X_PD NGD2VER_PD_9882 (.O (GTS) );
  endmodule
